# Created by MC2 : Version 2012.02.00.d on 2025/06/20, 22:37:44

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpuhddpsram_2012.02.00.d.170a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile 1P10M HKMG CU_ELK 0.9V				*/
# Memory Type    : TSMC 28nm High Performance Compact Mobile Ultra High Density Dual Port SRAM with d127 bit cell SVT Periphery */
# Library Name   : tsdn28hpcpuhdb32x16m4mwa (user specify : TSDN28HPCPUHDB32X16M4MWA)				*/
# Library Version: 170a												*/
# Generated Time : 2025/06/20, 22:37:43										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TSDN28HPCPUHDB32X16M4MWA
	CLASS BLOCK ;
	FOREIGN TSDN28HPCPUHDB32X16M4MWA 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 47.785 BY 57.850 ;
	SYMMETRY X Y ;
	PIN AA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 29.565 47.785 29.715 ;
			LAYER M2 ;
			RECT 47.605 29.565 47.785 29.715 ;
			LAYER M3 ;
			RECT 47.605 29.565 47.785 29.715 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[0]

	PIN AA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 32.115 47.785 32.265 ;
			LAYER M2 ;
			RECT 47.605 32.115 47.785 32.265 ;
			LAYER M1 ;
			RECT 47.605 32.115 47.785 32.265 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[1]

	PIN AA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 22.015 47.785 22.165 ;
			LAYER M3 ;
			RECT 47.605 22.015 47.785 22.165 ;
			LAYER M2 ;
			RECT 47.605 22.015 47.785 22.165 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[2]

	PIN AA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 23.465 47.785 23.615 ;
			LAYER M1 ;
			RECT 47.605 23.465 47.785 23.615 ;
			LAYER M3 ;
			RECT 47.605 23.465 47.785 23.615 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[3]

	PIN AA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 23.825 47.785 23.975 ;
			LAYER M2 ;
			RECT 47.605 23.825 47.785 23.975 ;
			LAYER M3 ;
			RECT 47.605 23.825 47.785 23.975 ;
		END
		ANTENNAGATEAREA 0.076800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.534300 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.076800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.845700 LAYER M2 ;
		ANTENNAMAXAREACAR 23.321800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.677200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.076800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.774000 LAYER M3 ;
		ANTENNAMAXAREACAR 27.573000 LAYER M3 ;
	END AA[4]

	PIN AB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 29.895 47.785 30.045 ;
			LAYER M3 ;
			RECT 47.605 29.895 47.785 30.045 ;
			LAYER M1 ;
			RECT 47.605 29.895 47.785 30.045 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[0]

	PIN AB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 31.785 47.785 31.935 ;
			LAYER M3 ;
			RECT 47.605 31.785 47.785 31.935 ;
			LAYER M1 ;
			RECT 47.605 31.785 47.785 31.935 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[1]

	PIN AB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 22.345 47.785 22.495 ;
			LAYER M3 ;
			RECT 47.605 22.345 47.785 22.495 ;
			LAYER M2 ;
			RECT 47.605 22.345 47.785 22.495 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[2]

	PIN AB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 23.135 47.785 23.285 ;
			LAYER M3 ;
			RECT 47.605 23.135 47.785 23.285 ;
			LAYER M2 ;
			RECT 47.605 23.135 47.785 23.285 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[3]

	PIN AB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 24.155 47.785 24.305 ;
			LAYER M2 ;
			RECT 47.605 24.155 47.785 24.305 ;
			LAYER M1 ;
			RECT 47.605 24.155 47.785 24.305 ;
		END
		ANTENNAGATEAREA 0.060300 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.437200 LAYER M1 ;
		ANTENNAMAXAREACAR 2.215600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.060300 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.812900 LAYER M2 ;
		ANTENNAMAXAREACAR 34.966700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.866700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.060300 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.869800 LAYER M3 ;
		ANTENNAMAXAREACAR 47.190400 LAYER M3 ;
	END AB[4]

	PIN AWT
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 47.230 47.785 47.380 ;
			LAYER M2 ;
			RECT 47.605 47.230 47.785 47.380 ;
			LAYER M1 ;
			RECT 47.605 47.230 47.785 47.380 ;
		END
		ANTENNAGATEAREA 0.129000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.279100 LAYER M1 ;
		ANTENNAMAXAREACAR 0.723600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.151200 LAYER VIA1 ;
		ANTENNAGATEAREA 0.129000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.591000 LAYER M2 ;
		ANTENNAMAXAREACAR 5.305000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.201600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.129000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.514300 LAYER M3 ;
	END AWT

	PIN BWEBA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 1.525 47.785 1.675 ;
			LAYER M2 ;
			RECT 47.605 1.525 47.785 1.675 ;
			LAYER M3 ;
			RECT 47.605 1.525 47.785 1.675 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[0]

	PIN BWEBA[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 42.940 47.785 43.090 ;
			LAYER M1 ;
			RECT 47.605 42.940 47.785 43.090 ;
			LAYER M2 ;
			RECT 47.605 42.940 47.785 43.090 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[10]

	PIN BWEBA[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 45.910 47.785 46.060 ;
			LAYER M3 ;
			RECT 47.605 45.910 47.785 46.060 ;
			LAYER M1 ;
			RECT 47.605 45.910 47.785 46.060 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[11]

	PIN BWEBA[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 48.220 47.785 48.370 ;
			LAYER M2 ;
			RECT 47.605 48.220 47.785 48.370 ;
			LAYER M1 ;
			RECT 47.605 48.220 47.785 48.370 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[12]

	PIN BWEBA[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 50.205 47.785 50.355 ;
			LAYER M3 ;
			RECT 47.605 50.205 47.785 50.355 ;
			LAYER M1 ;
			RECT 47.605 50.205 47.785 50.355 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[13]

	PIN BWEBA[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 52.525 47.785 52.675 ;
			LAYER M2 ;
			RECT 47.605 52.525 47.785 52.675 ;
			LAYER M3 ;
			RECT 47.605 52.525 47.785 52.675 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[14]

	PIN BWEBA[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 54.845 47.785 54.995 ;
			LAYER M1 ;
			RECT 47.605 54.845 47.785 54.995 ;
			LAYER M2 ;
			RECT 47.605 54.845 47.785 54.995 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[15]

	PIN BWEBA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 3.845 47.785 3.995 ;
			LAYER M3 ;
			RECT 47.605 3.845 47.785 3.995 ;
			LAYER M1 ;
			RECT 47.605 3.845 47.785 3.995 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[1]

	PIN BWEBA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 6.165 47.785 6.315 ;
			LAYER M2 ;
			RECT 47.605 6.165 47.785 6.315 ;
			LAYER M1 ;
			RECT 47.605 6.165 47.785 6.315 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[2]

	PIN BWEBA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 8.485 47.785 8.635 ;
			LAYER M3 ;
			RECT 47.605 8.485 47.785 8.635 ;
			LAYER M1 ;
			RECT 47.605 8.485 47.785 8.635 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[3]

	PIN BWEBA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 10.795 47.785 10.945 ;
			LAYER M1 ;
			RECT 47.605 10.795 47.785 10.945 ;
			LAYER M2 ;
			RECT 47.605 10.795 47.785 10.945 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[4]

	PIN BWEBA[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 12.775 47.785 12.925 ;
			LAYER M2 ;
			RECT 47.605 12.775 47.785 12.925 ;
			LAYER M3 ;
			RECT 47.605 12.775 47.785 12.925 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[5]

	PIN BWEBA[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 15.670 47.785 15.820 ;
			LAYER M2 ;
			RECT 47.605 15.670 47.785 15.820 ;
			LAYER M1 ;
			RECT 47.605 15.670 47.785 15.820 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[6]

	PIN BWEBA[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 17.670 47.785 17.820 ;
			LAYER M1 ;
			RECT 47.605 17.670 47.785 17.820 ;
			LAYER M2 ;
			RECT 47.605 17.670 47.785 17.820 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[7]

	PIN BWEBA[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 38.020 47.785 38.170 ;
			LAYER M2 ;
			RECT 47.605 38.020 47.785 38.170 ;
			LAYER M1 ;
			RECT 47.605 38.020 47.785 38.170 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[8]

	PIN BWEBA[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 40.630 47.785 40.780 ;
			LAYER M2 ;
			RECT 47.605 40.630 47.785 40.780 ;
			LAYER M3 ;
			RECT 47.605 40.630 47.785 40.780 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.177600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.776000 LAYER M2 ;
		ANTENNAMAXAREACAR 73.370400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.242700 LAYER M3 ;
		ANTENNAMAXAREACAR 75.870400 LAYER M3 ;
	END BWEBA[9]

	PIN BWEBB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 1.195 47.785 1.345 ;
			LAYER M1 ;
			RECT 47.605 1.195 47.785 1.345 ;
			LAYER M2 ;
			RECT 47.605 1.195 47.785 1.345 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[0]

	PIN BWEBB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 42.610 47.785 42.760 ;
			LAYER M1 ;
			RECT 47.605 42.610 47.785 42.760 ;
			LAYER M3 ;
			RECT 47.605 42.610 47.785 42.760 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[10]

	PIN BWEBB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 45.580 47.785 45.730 ;
			LAYER M2 ;
			RECT 47.605 45.580 47.785 45.730 ;
			LAYER M1 ;
			RECT 47.605 45.580 47.785 45.730 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[11]

	PIN BWEBB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 47.890 47.785 48.040 ;
			LAYER M2 ;
			RECT 47.605 47.890 47.785 48.040 ;
			LAYER M3 ;
			RECT 47.605 47.890 47.785 48.040 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[12]

	PIN BWEBB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 49.875 47.785 50.025 ;
			LAYER M2 ;
			RECT 47.605 49.875 47.785 50.025 ;
			LAYER M1 ;
			RECT 47.605 49.875 47.785 50.025 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[13]

	PIN BWEBB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 52.195 47.785 52.345 ;
			LAYER M3 ;
			RECT 47.605 52.195 47.785 52.345 ;
			LAYER M2 ;
			RECT 47.605 52.195 47.785 52.345 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[14]

	PIN BWEBB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 54.515 47.785 54.665 ;
			LAYER M3 ;
			RECT 47.605 54.515 47.785 54.665 ;
			LAYER M2 ;
			RECT 47.605 54.515 47.785 54.665 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[15]

	PIN BWEBB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 3.515 47.785 3.665 ;
			LAYER M3 ;
			RECT 47.605 3.515 47.785 3.665 ;
			LAYER M1 ;
			RECT 47.605 3.515 47.785 3.665 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[1]

	PIN BWEBB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 5.835 47.785 5.985 ;
			LAYER M1 ;
			RECT 47.605 5.835 47.785 5.985 ;
			LAYER M2 ;
			RECT 47.605 5.835 47.785 5.985 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[2]

	PIN BWEBB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 8.155 47.785 8.305 ;
			LAYER M1 ;
			RECT 47.605 8.155 47.785 8.305 ;
			LAYER M3 ;
			RECT 47.605 8.155 47.785 8.305 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[3]

	PIN BWEBB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 10.465 47.785 10.615 ;
			LAYER M1 ;
			RECT 47.605 10.465 47.785 10.615 ;
			LAYER M2 ;
			RECT 47.605 10.465 47.785 10.615 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[4]

	PIN BWEBB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 12.445 47.785 12.595 ;
			LAYER M3 ;
			RECT 47.605 12.445 47.785 12.595 ;
			LAYER M2 ;
			RECT 47.605 12.445 47.785 12.595 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[5]

	PIN BWEBB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 15.340 47.785 15.490 ;
			LAYER M2 ;
			RECT 47.605 15.340 47.785 15.490 ;
			LAYER M3 ;
			RECT 47.605 15.340 47.785 15.490 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[6]

	PIN BWEBB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 17.320 47.785 17.470 ;
			LAYER M3 ;
			RECT 47.605 17.320 47.785 17.470 ;
			LAYER M2 ;
			RECT 47.605 17.320 47.785 17.470 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[7]

	PIN BWEBB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 37.690 47.785 37.840 ;
			LAYER M1 ;
			RECT 47.605 37.690 47.785 37.840 ;
			LAYER M3 ;
			RECT 47.605 37.690 47.785 37.840 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[8]

	PIN BWEBB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 40.300 47.785 40.450 ;
			LAYER M3 ;
			RECT 47.605 40.300 47.785 40.450 ;
			LAYER M1 ;
			RECT 47.605 40.300 47.785 40.450 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.349700 LAYER M1 ;
		ANTENNAMAXAREACAR 19.050900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.829000 LAYER M2 ;
		ANTENNAMAXAREACAR 90.180600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.187500 LAYER M3 ;
		ANTENNAMAXAREACAR 92.680600 LAYER M3 ;
	END BWEBB[9]

	PIN CEBA
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 36.700 47.785 36.850 ;
			LAYER M3 ;
			RECT 47.605 36.700 47.785 36.850 ;
			LAYER M1 ;
			RECT 47.605 36.700 47.785 36.850 ;
		END
		ANTENNAGATEAREA 0.068100 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.266600 LAYER M1 ;
		ANTENNAMAXAREACAR 2.847400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.223400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.068100 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.577800 LAYER M2 ;
		ANTENNAMAXAREACAR 10.714500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.318800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.068100 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.261500 LAYER M3 ;
		ANTENNAMAXAREACAR 12.155100 LAYER M3 ;
	END CEBA

	PIN CEBB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 37.030 47.785 37.180 ;
			LAYER M1 ;
			RECT 47.605 37.030 47.785 37.180 ;
			LAYER M3 ;
			RECT 47.605 37.030 47.785 37.180 ;
		END
		ANTENNAGATEAREA 0.029100 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.342200 LAYER M1 ;
		ANTENNAMAXAREACAR 10.096200 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.223400 LAYER VIA1 ;
		ANTENNAGATEAREA 0.029100 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.644400 LAYER M2 ;
		ANTENNAMAXAREACAR 32.239700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.446700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.029100 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 33.167500 LAYER M3 ;
	END CEBB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 34.720 47.785 34.870 ;
			LAYER M1 ;
			RECT 47.605 34.720 47.785 34.870 ;
			LAYER M3 ;
			RECT 47.605 34.720 47.785 34.870 ;
		END
		ANTENNAGATEAREA 0.394500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.757100 LAYER M1 ;
		ANTENNAMAXAREACAR 3.389600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.656600 LAYER VIA1 ;
		ANTENNAGATEAREA 0.394500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.828600 LAYER M2 ;
		ANTENNAMAXAREACAR 8.667400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.039000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.313100 LAYER VIA2 ;
		ANTENNAGATEAREA 0.394500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.952600 LAYER M3 ;
		ANTENNAMAXAREACAR 11.082000 LAYER M3 ;
	END CLK

	PIN DA[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 2.855 47.785 3.005 ;
			LAYER M2 ;
			RECT 47.605 2.855 47.785 3.005 ;
			LAYER M3 ;
			RECT 47.605 2.855 47.785 3.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[0]

	PIN DA[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 44.920 47.785 45.070 ;
			LAYER M3 ;
			RECT 47.605 44.920 47.785 45.070 ;
			LAYER M1 ;
			RECT 47.605 44.920 47.785 45.070 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[10]

	PIN DA[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 46.900 47.785 47.050 ;
			LAYER M3 ;
			RECT 47.605 46.900 47.785 47.050 ;
			LAYER M1 ;
			RECT 47.605 46.900 47.785 47.050 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[11]

	PIN DA[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 49.215 47.785 49.365 ;
			LAYER M3 ;
			RECT 47.605 49.215 47.785 49.365 ;
			LAYER M2 ;
			RECT 47.605 49.215 47.785 49.365 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[12]

	PIN DA[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 51.535 47.785 51.685 ;
			LAYER M2 ;
			RECT 47.605 51.535 47.785 51.685 ;
			LAYER M3 ;
			RECT 47.605 51.535 47.785 51.685 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[13]

	PIN DA[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 53.855 47.785 54.005 ;
			LAYER M2 ;
			RECT 47.605 53.855 47.785 54.005 ;
			LAYER M3 ;
			RECT 47.605 53.855 47.785 54.005 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[14]

	PIN DA[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 56.175 47.785 56.325 ;
			LAYER M1 ;
			RECT 47.605 56.175 47.785 56.325 ;
			LAYER M2 ;
			RECT 47.605 56.175 47.785 56.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[15]

	PIN DA[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 5.175 47.785 5.325 ;
			LAYER M3 ;
			RECT 47.605 5.175 47.785 5.325 ;
			LAYER M1 ;
			RECT 47.605 5.175 47.785 5.325 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[1]

	PIN DA[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 7.495 47.785 7.645 ;
			LAYER M1 ;
			RECT 47.605 7.495 47.785 7.645 ;
			LAYER M2 ;
			RECT 47.605 7.495 47.785 7.645 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[2]

	PIN DA[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 9.475 47.785 9.625 ;
			LAYER M3 ;
			RECT 47.605 9.475 47.785 9.625 ;
			LAYER M2 ;
			RECT 47.605 9.475 47.785 9.625 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[3]

	PIN DA[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 11.785 47.785 11.935 ;
			LAYER M3 ;
			RECT 47.605 11.785 47.785 11.935 ;
			LAYER M1 ;
			RECT 47.605 11.785 47.785 11.935 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[4]

	PIN DA[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 13.765 47.785 13.915 ;
			LAYER M3 ;
			RECT 47.605 13.765 47.785 13.915 ;
			LAYER M2 ;
			RECT 47.605 13.765 47.785 13.915 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[5]

	PIN DA[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 16.660 47.785 16.810 ;
			LAYER M1 ;
			RECT 47.605 16.660 47.785 16.810 ;
			LAYER M2 ;
			RECT 47.605 16.660 47.785 16.810 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[6]

	PIN DA[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 18.705 47.785 18.855 ;
			LAYER M2 ;
			RECT 47.605 18.705 47.785 18.855 ;
			LAYER M3 ;
			RECT 47.605 18.705 47.785 18.855 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[7]

	PIN DA[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 39.010 47.785 39.160 ;
			LAYER M1 ;
			RECT 47.605 39.010 47.785 39.160 ;
			LAYER M2 ;
			RECT 47.605 39.010 47.785 39.160 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[8]

	PIN DA[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 41.620 47.785 41.770 ;
			LAYER M1 ;
			RECT 47.605 41.620 47.785 41.770 ;
			LAYER M3 ;
			RECT 47.605 41.620 47.785 41.770 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.131300 LAYER M1 ;
		ANTENNAMAXAREACAR 2.398100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.601900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.868500 LAYER M2 ;
		ANTENNAMAXAREACAR 82.814800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.220000 LAYER M3 ;
		ANTENNAMAXAREACAR 85.314800 LAYER M3 ;
	END DA[9]

	PIN DB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 3.185 47.785 3.335 ;
			LAYER M1 ;
			RECT 47.605 3.185 47.785 3.335 ;
			LAYER M2 ;
			RECT 47.605 3.185 47.785 3.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[0]

	PIN DB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 45.250 47.785 45.400 ;
			LAYER M1 ;
			RECT 47.605 45.250 47.785 45.400 ;
			LAYER M3 ;
			RECT 47.605 45.250 47.785 45.400 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[10]

	PIN DB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 47.560 47.785 47.710 ;
			LAYER M3 ;
			RECT 47.605 47.560 47.785 47.710 ;
			LAYER M2 ;
			RECT 47.605 47.560 47.785 47.710 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[11]

	PIN DB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 49.545 47.785 49.695 ;
			LAYER M2 ;
			RECT 47.605 49.545 47.785 49.695 ;
			LAYER M3 ;
			RECT 47.605 49.545 47.785 49.695 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[12]

	PIN DB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 51.865 47.785 52.015 ;
			LAYER M3 ;
			RECT 47.605 51.865 47.785 52.015 ;
			LAYER M1 ;
			RECT 47.605 51.865 47.785 52.015 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[13]

	PIN DB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 54.185 47.785 54.335 ;
			LAYER M2 ;
			RECT 47.605 54.185 47.785 54.335 ;
			LAYER M1 ;
			RECT 47.605 54.185 47.785 54.335 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[14]

	PIN DB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 56.505 47.785 56.655 ;
			LAYER M1 ;
			RECT 47.605 56.505 47.785 56.655 ;
			LAYER M2 ;
			RECT 47.605 56.505 47.785 56.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[15]

	PIN DB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 5.505 47.785 5.655 ;
			LAYER M1 ;
			RECT 47.605 5.505 47.785 5.655 ;
			LAYER M2 ;
			RECT 47.605 5.505 47.785 5.655 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[1]

	PIN DB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 7.825 47.785 7.975 ;
			LAYER M1 ;
			RECT 47.605 7.825 47.785 7.975 ;
			LAYER M2 ;
			RECT 47.605 7.825 47.785 7.975 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[2]

	PIN DB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 10.135 47.785 10.285 ;
			LAYER M2 ;
			RECT 47.605 10.135 47.785 10.285 ;
			LAYER M1 ;
			RECT 47.605 10.135 47.785 10.285 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[3]

	PIN DB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 12.115 47.785 12.265 ;
			LAYER M1 ;
			RECT 47.605 12.115 47.785 12.265 ;
			LAYER M3 ;
			RECT 47.605 12.115 47.785 12.265 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[4]

	PIN DB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 15.010 47.785 15.160 ;
			LAYER M3 ;
			RECT 47.605 15.010 47.785 15.160 ;
			LAYER M2 ;
			RECT 47.605 15.010 47.785 15.160 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[5]

	PIN DB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 16.990 47.785 17.140 ;
			LAYER M1 ;
			RECT 47.605 16.990 47.785 17.140 ;
			LAYER M3 ;
			RECT 47.605 16.990 47.785 17.140 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[6]

	PIN DB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 19.035 47.785 19.185 ;
			LAYER M3 ;
			RECT 47.605 19.035 47.785 19.185 ;
			LAYER M1 ;
			RECT 47.605 19.035 47.785 19.185 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[7]

	PIN DB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 39.970 47.785 40.120 ;
			LAYER M3 ;
			RECT 47.605 39.970 47.785 40.120 ;
			LAYER M1 ;
			RECT 47.605 39.970 47.785 40.120 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[8]

	PIN DB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 42.280 47.785 42.430 ;
			LAYER M3 ;
			RECT 47.605 42.280 47.785 42.430 ;
			LAYER M1 ;
			RECT 47.605 42.280 47.785 42.430 ;
		END
		ANTENNAGATEAREA 0.010800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.344500 LAYER M1 ;
		ANTENNAMAXAREACAR 18.476900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 1.203700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.010800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.875900 LAYER M2 ;
		ANTENNAMAXAREACAR 89.032400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.805600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.010800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.129300 LAYER M3 ;
		ANTENNAMAXAREACAR 91.532400 LAYER M3 ;
	END DB[9]

	PIN PTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 34.060 47.785 34.210 ;
			LAYER M3 ;
			RECT 47.605 34.060 47.785 34.210 ;
			LAYER M1 ;
			RECT 47.605 34.060 47.785 34.210 ;
		END
		ANTENNAGATEAREA 0.015900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.219900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.012600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.408800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.015900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483500 LAYER M2 ;
		ANTENNAMAXAREACAR 31.421400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.817600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.015900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121200 LAYER M3 ;
		ANTENNAMAXAREACAR 33.119500 LAYER M3 ;
	END PTSEL[0]

	PIN PTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 34.390 47.785 34.540 ;
			LAYER M3 ;
			RECT 47.605 34.390 47.785 34.540 ;
			LAYER M1 ;
			RECT 47.605 34.390 47.785 34.540 ;
		END
		ANTENNAGATEAREA 0.015900 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.219900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.012600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.408800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.015900 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.483500 LAYER M2 ;
		ANTENNAMAXAREACAR 31.421400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.817600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.015900 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.121200 LAYER M3 ;
		ANTENNAMAXAREACAR 33.119500 LAYER M3 ;
	END PTSEL[1]

	PIN QA[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 1.860 47.785 2.010 ;
			LAYER M3 ;
			RECT 47.605 1.860 47.785 2.010 ;
			LAYER M1 ;
			RECT 47.605 1.860 47.785 2.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[0]

	PIN QA[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 43.270 47.785 43.420 ;
			LAYER M1 ;
			RECT 47.605 43.270 47.785 43.420 ;
			LAYER M2 ;
			RECT 47.605 43.270 47.785 43.420 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[10]

	PIN QA[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 46.240 47.785 46.390 ;
			LAYER M1 ;
			RECT 47.605 46.240 47.785 46.390 ;
			LAYER M2 ;
			RECT 47.605 46.240 47.785 46.390 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[11]

	PIN QA[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 48.550 47.785 48.700 ;
			LAYER M1 ;
			RECT 47.605 48.550 47.785 48.700 ;
			LAYER M2 ;
			RECT 47.605 48.550 47.785 48.700 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[12]

	PIN QA[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 50.540 47.785 50.690 ;
			LAYER M3 ;
			RECT 47.605 50.540 47.785 50.690 ;
			LAYER M1 ;
			RECT 47.605 50.540 47.785 50.690 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[13]

	PIN QA[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 52.860 47.785 53.010 ;
			LAYER M1 ;
			RECT 47.605 52.860 47.785 53.010 ;
			LAYER M3 ;
			RECT 47.605 52.860 47.785 53.010 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[14]

	PIN QA[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 55.180 47.785 55.330 ;
			LAYER M3 ;
			RECT 47.605 55.180 47.785 55.330 ;
			LAYER M1 ;
			RECT 47.605 55.180 47.785 55.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[15]

	PIN QA[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 4.180 47.785 4.330 ;
			LAYER M1 ;
			RECT 47.605 4.180 47.785 4.330 ;
			LAYER M2 ;
			RECT 47.605 4.180 47.785 4.330 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[1]

	PIN QA[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 6.500 47.785 6.650 ;
			LAYER M1 ;
			RECT 47.605 6.500 47.785 6.650 ;
			LAYER M2 ;
			RECT 47.605 6.500 47.785 6.650 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[2]

	PIN QA[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 8.815 47.785 8.965 ;
			LAYER M3 ;
			RECT 47.605 8.815 47.785 8.965 ;
			LAYER M1 ;
			RECT 47.605 8.815 47.785 8.965 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[3]

	PIN QA[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 11.125 47.785 11.275 ;
			LAYER M2 ;
			RECT 47.605 11.125 47.785 11.275 ;
			LAYER M3 ;
			RECT 47.605 11.125 47.785 11.275 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[4]

	PIN QA[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 13.105 47.785 13.255 ;
			LAYER M1 ;
			RECT 47.605 13.105 47.785 13.255 ;
			LAYER M2 ;
			RECT 47.605 13.105 47.785 13.255 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[5]

	PIN QA[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 16.000 47.785 16.150 ;
			LAYER M2 ;
			RECT 47.605 16.000 47.785 16.150 ;
			LAYER M1 ;
			RECT 47.605 16.000 47.785 16.150 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[6]

	PIN QA[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 18.000 47.785 18.150 ;
			LAYER M1 ;
			RECT 47.605 18.000 47.785 18.150 ;
			LAYER M3 ;
			RECT 47.605 18.000 47.785 18.150 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[7]

	PIN QA[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 38.350 47.785 38.500 ;
			LAYER M1 ;
			RECT 47.605 38.350 47.785 38.500 ;
			LAYER M3 ;
			RECT 47.605 38.350 47.785 38.500 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[8]

	PIN QA[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 40.960 47.785 41.110 ;
			LAYER M1 ;
			RECT 47.605 40.960 47.785 41.110 ;
			LAYER M2 ;
			RECT 47.605 40.960 47.785 41.110 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.272700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.901600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.239100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.641200 LAYER M4 ;
	END QA[9]

	PIN QB[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 2.525 47.785 2.675 ;
			LAYER M1 ;
			RECT 47.605 2.525 47.785 2.675 ;
			LAYER M3 ;
			RECT 47.605 2.525 47.785 2.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[0]

	PIN QB[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 44.590 47.785 44.740 ;
			LAYER M3 ;
			RECT 47.605 44.590 47.785 44.740 ;
			LAYER M1 ;
			RECT 47.605 44.590 47.785 44.740 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[10]

	PIN QB[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 46.570 47.785 46.720 ;
			LAYER M2 ;
			RECT 47.605 46.570 47.785 46.720 ;
			LAYER M3 ;
			RECT 47.605 46.570 47.785 46.720 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[11]

	PIN QB[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 48.885 47.785 49.035 ;
			LAYER M3 ;
			RECT 47.605 48.885 47.785 49.035 ;
			LAYER M1 ;
			RECT 47.605 48.885 47.785 49.035 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[12]

	PIN QB[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 51.205 47.785 51.355 ;
			LAYER M1 ;
			RECT 47.605 51.205 47.785 51.355 ;
			LAYER M2 ;
			RECT 47.605 51.205 47.785 51.355 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[13]

	PIN QB[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 53.525 47.785 53.675 ;
			LAYER M1 ;
			RECT 47.605 53.525 47.785 53.675 ;
			LAYER M2 ;
			RECT 47.605 53.525 47.785 53.675 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[14]

	PIN QB[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 55.845 47.785 55.995 ;
			LAYER M2 ;
			RECT 47.605 55.845 47.785 55.995 ;
			LAYER M1 ;
			RECT 47.605 55.845 47.785 55.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[15]

	PIN QB[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 4.845 47.785 4.995 ;
			LAYER M1 ;
			RECT 47.605 4.845 47.785 4.995 ;
			LAYER M2 ;
			RECT 47.605 4.845 47.785 4.995 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[1]

	PIN QB[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 7.165 47.785 7.315 ;
			LAYER M1 ;
			RECT 47.605 7.165 47.785 7.315 ;
			LAYER M2 ;
			RECT 47.605 7.165 47.785 7.315 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[2]

	PIN QB[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 9.145 47.785 9.295 ;
			LAYER M1 ;
			RECT 47.605 9.145 47.785 9.295 ;
			LAYER M3 ;
			RECT 47.605 9.145 47.785 9.295 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[3]

	PIN QB[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 11.455 47.785 11.605 ;
			LAYER M1 ;
			RECT 47.605 11.455 47.785 11.605 ;
			LAYER M2 ;
			RECT 47.605 11.455 47.785 11.605 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[4]

	PIN QB[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 13.435 47.785 13.585 ;
			LAYER M1 ;
			RECT 47.605 13.435 47.785 13.585 ;
			LAYER M3 ;
			RECT 47.605 13.435 47.785 13.585 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[5]

	PIN QB[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 16.330 47.785 16.480 ;
			LAYER M2 ;
			RECT 47.605 16.330 47.785 16.480 ;
			LAYER M1 ;
			RECT 47.605 16.330 47.785 16.480 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[6]

	PIN QB[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 18.375 47.785 18.525 ;
			LAYER M2 ;
			RECT 47.605 18.375 47.785 18.525 ;
			LAYER M3 ;
			RECT 47.605 18.375 47.785 18.525 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[7]

	PIN QB[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 38.680 47.785 38.830 ;
			LAYER M3 ;
			RECT 47.605 38.680 47.785 38.830 ;
			LAYER M1 ;
			RECT 47.605 38.680 47.785 38.830 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[8]

	PIN QB[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 41.290 47.785 41.440 ;
			LAYER M2 ;
			RECT 47.605 41.290 47.785 41.440 ;
			LAYER M1 ;
			RECT 47.605 41.290 47.785 41.440 ;
		END
		ANTENNADIFFAREA 0.155000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.173700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNADIFFAREA 0.155000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.000500 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.058500 LAYER VIA2 ;
		ANTENNADIFFAREA 0.155000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.443500 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA3 ;
		ANTENNADIFFAREA 0.155000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 0.642900 LAYER M4 ;
	END QB[9]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 43.930 47.785 44.080 ;
			LAYER M2 ;
			RECT 47.605 43.930 47.785 44.080 ;
			LAYER M1 ;
			RECT 47.605 43.930 47.785 44.080 ;
		END
		ANTENNAGATEAREA 0.045600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.275900 LAYER M1 ;
		ANTENNAMAXAREACAR 7.227300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.393900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.045600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.199800 LAYER M2 ;
		ANTENNAMAXAREACAR 11.181800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.787900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.045600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.090400 LAYER M3 ;
		ANTENNAMAXAREACAR 12.818200 LAYER M3 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 44.260 47.785 44.410 ;
			LAYER M2 ;
			RECT 47.605 44.260 47.785 44.410 ;
			LAYER M3 ;
			RECT 47.605 44.260 47.785 44.410 ;
		END
		ANTENNAGATEAREA 0.045600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.275900 LAYER M1 ;
		ANTENNAMAXAREACAR 7.227300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.393900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.045600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.199800 LAYER M2 ;
		ANTENNAMAXAREACAR 11.181800 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.787900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.045600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.090400 LAYER M3 ;
		ANTENNAMAXAREACAR 12.818200 LAYER M3 ;
	END RTSEL[1]

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 1.395 47.395 1.725 ;
			LAYER M4 ;
			RECT 0.000 3.715 47.395 4.045 ;
			LAYER M4 ;
			RECT 0.000 6.035 47.395 6.365 ;
			LAYER M4 ;
			RECT 0.000 8.355 47.395 8.685 ;
			LAYER M4 ;
			RECT 0.000 10.675 47.395 11.005 ;
			LAYER M4 ;
			RECT 0.000 12.995 47.395 13.325 ;
			LAYER M4 ;
			RECT 0.000 15.315 47.395 15.645 ;
			LAYER M4 ;
			RECT 0.000 17.635 47.395 17.965 ;
			LAYER M4 ;
			RECT 0.000 19.985 47.395 20.290 ;
			LAYER M4 ;
			RECT 0.000 23.850 47.395 24.400 ;
			LAYER M4 ;
			RECT 0.000 24.905 47.395 25.325 ;
			LAYER M4 ;
			RECT 0.000 26.870 47.395 27.440 ;
			LAYER M4 ;
			RECT 0.000 27.570 47.395 28.140 ;
			LAYER M4 ;
			RECT 24.150 30.280 47.395 30.930 ;
			LAYER M4 ;
			RECT 0.000 32.030 47.395 32.680 ;
			LAYER M4 ;
			RECT 0.000 34.825 47.395 35.475 ;
			LAYER M4 ;
			RECT 0.000 35.625 47.395 35.935 ;
			LAYER M4 ;
			RECT 0.000 38.475 47.395 38.805 ;
			LAYER M4 ;
			RECT 0.000 40.795 47.395 41.125 ;
			LAYER M4 ;
			RECT 0.000 43.115 47.395 43.445 ;
			LAYER M4 ;
			RECT 0.000 45.435 47.395 45.765 ;
			LAYER M4 ;
			RECT 0.000 47.755 47.395 48.085 ;
			LAYER M4 ;
			RECT 0.000 50.075 47.395 50.405 ;
			LAYER M4 ;
			RECT 0.000 52.395 47.395 52.725 ;
			LAYER M4 ;
			RECT 0.000 54.715 47.395 55.045 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 2.805 47.395 3.185 ;
			LAYER M4 ;
			RECT 0.000 5.125 47.395 5.505 ;
			LAYER M4 ;
			RECT 0.000 7.445 47.395 7.825 ;
			LAYER M4 ;
			RECT 0.000 9.765 47.395 10.145 ;
			LAYER M4 ;
			RECT 0.000 12.085 47.395 12.465 ;
			LAYER M4 ;
			RECT 0.000 14.405 47.395 14.785 ;
			LAYER M4 ;
			RECT 0.000 16.725 47.395 17.105 ;
			LAYER M4 ;
			RECT 0.000 19.045 47.395 19.425 ;
			LAYER M4 ;
			RECT 21.525 22.310 47.395 23.090 ;
			LAYER M4 ;
			RECT 0.000 25.470 47.395 26.040 ;
			LAYER M4 ;
			RECT 0.000 26.170 47.395 26.740 ;
			LAYER M4 ;
			RECT 0.000 28.400 47.395 29.050 ;
			LAYER M4 ;
			RECT 24.150 29.480 47.395 30.130 ;
			LAYER M4 ;
			RECT 0.000 31.310 47.395 31.880 ;
			LAYER M4 ;
			RECT 0.000 39.885 47.395 40.265 ;
			LAYER M4 ;
			RECT 0.000 42.205 47.395 42.585 ;
			LAYER M4 ;
			RECT 0.000 44.525 47.395 44.905 ;
			LAYER M4 ;
			RECT 0.000 46.845 47.395 47.225 ;
			LAYER M4 ;
			RECT 0.000 49.165 47.395 49.545 ;
			LAYER M4 ;
			RECT 0.000 51.485 47.395 51.865 ;
			LAYER M4 ;
			RECT 0.000 53.805 47.395 54.185 ;
			LAYER M4 ;
			RECT 0.000 56.125 47.395 56.505 ;
		END
	END VSS

	PIN WEBA
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 32.445 47.785 32.595 ;
			LAYER M1 ;
			RECT 47.605 32.445 47.785 32.595 ;
			LAYER M2 ;
			RECT 47.605 32.445 47.785 32.595 ;
		END
		ANTENNAGATEAREA 0.039000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.170000 LAYER M1 ;
		ANTENNAMAXAREACAR 3.116700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.166700 LAYER VIA1 ;
		ANTENNAGATEAREA 0.039000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.530800 LAYER M2 ;
		ANTENNAMAXAREACAR 15.783300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.333300 LAYER VIA2 ;
		ANTENNAGATEAREA 0.039000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.122900 LAYER M3 ;
		ANTENNAMAXAREACAR 17.051300 LAYER M3 ;
	END WEBA

	PIN WEBB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 47.605 32.775 47.785 32.925 ;
			LAYER M1 ;
			RECT 47.605 32.775 47.785 32.925 ;
			LAYER M2 ;
			RECT 47.605 32.775 47.785 32.925 ;
		END
		ANTENNAGATEAREA 0.022500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.088700 LAYER M1 ;
		ANTENNAMAXAREACAR 1.788900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.288900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.022500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.465500 LAYER M2 ;
		ANTENNAMAXAREACAR 20.633300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.577800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.022500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.080200 LAYER M3 ;
		ANTENNAMAXAREACAR 21.833300 LAYER M3 ;
	END WEBB

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 47.605 37.355 47.785 37.505 ;
			LAYER M2 ;
			RECT 47.605 37.355 47.785 37.505 ;
			LAYER M3 ;
			RECT 47.605 37.355 47.785 37.505 ;
		END
		ANTENNAGATEAREA 0.022500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.073500 LAYER M1 ;
		ANTENNAMAXAREACAR 1.111100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.288900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.022500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.383200 LAYER M2 ;
		ANTENNAMAXAREACAR 17.766700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.577800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.022500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.202700 LAYER M3 ;
		ANTENNAMAXAREACAR 18.966700 LAYER M3 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.605 36.370 47.785 36.520 ;
			LAYER M1 ;
			RECT 47.605 36.370 47.785 36.520 ;
			LAYER M3 ;
			RECT 47.605 36.370 47.785 36.520 ;
		END
		ANTENNAGATEAREA 0.022500 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.073500 LAYER M1 ;
		ANTENNAMAXAREACAR 1.111100 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.288900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.022500 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.383200 LAYER M2 ;
		ANTENNAMAXAREACAR 17.766700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.577800 LAYER VIA2 ;
		ANTENNAGATEAREA 0.022500 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.202700 LAYER M3 ;
		ANTENNAMAXAREACAR 18.966700 LAYER M3 ;
	END WTSEL[1]

	OBS
		# Promoted blockages
		LAYER M1 ;
		RECT 47.605 56.715 47.785 57.850 ;
		LAYER VIA3 ;
		RECT 47.605 56.735 47.785 57.850 ;
		LAYER VIA3 ;
		RECT 47.605 46.140 47.785 46.160 ;
		LAYER M2 ;
		RECT 47.605 54.745 47.785 54.765 ;
		LAYER M1 ;
		RECT 47.605 54.725 47.785 54.785 ;
		LAYER M3 ;
		RECT 47.605 46.140 47.785 46.160 ;
		LAYER M3 ;
		RECT 47.605 45.810 47.785 45.830 ;
		LAYER M1 ;
		RECT 47.605 46.120 47.785 46.180 ;
		LAYER M2 ;
		RECT 47.605 46.140 47.785 46.160 ;
		LAYER M1 ;
		RECT 47.605 45.790 47.785 45.850 ;
		LAYER M2 ;
		RECT 47.605 45.810 47.785 45.830 ;
		LAYER M2 ;
		RECT 47.605 45.150 47.785 45.170 ;
		LAYER VIA3 ;
		RECT 47.605 45.810 47.785 45.830 ;
		LAYER M3 ;
		RECT 47.605 45.150 47.785 45.170 ;
		LAYER VIA3 ;
		RECT 47.605 45.150 47.785 45.170 ;
		LAYER M3 ;
		RECT 47.605 56.405 47.785 56.425 ;
		LAYER M1 ;
		RECT 47.605 45.130 47.785 45.190 ;
		LAYER M1 ;
		RECT 47.605 44.800 47.785 44.860 ;
		LAYER M2 ;
		RECT 47.605 44.820 47.785 44.840 ;
		LAYER M3 ;
		RECT 47.605 44.820 47.785 44.840 ;
		LAYER VIA3 ;
		RECT 47.605 44.820 47.785 44.840 ;
		LAYER M2 ;
		RECT 47.605 45.480 47.785 45.500 ;
		LAYER M3 ;
		RECT 47.605 45.480 47.785 45.500 ;
		LAYER VIA3 ;
		RECT 47.605 45.480 47.785 45.500 ;
		LAYER M1 ;
		RECT 47.605 45.460 47.785 45.520 ;
		LAYER M1 ;
		RECT 47.605 49.095 47.785 49.155 ;
		LAYER VIA3 ;
		RECT 47.605 48.450 47.785 48.470 ;
		LAYER M3 ;
		RECT 47.605 48.450 47.785 48.470 ;
		LAYER M2 ;
		RECT 47.605 49.115 47.785 49.135 ;
		LAYER M3 ;
		RECT 47.605 49.115 47.785 49.135 ;
		LAYER VIA3 ;
		RECT 47.605 49.115 47.785 49.135 ;
		LAYER M2 ;
		RECT 47.605 48.780 47.785 48.805 ;
		LAYER VIA3 ;
		RECT 47.605 48.780 47.785 48.805 ;
		LAYER M3 ;
		RECT 47.605 48.780 47.785 48.805 ;
		LAYER M1 ;
		RECT 47.605 48.760 47.785 48.825 ;
		LAYER M3 ;
		RECT 47.605 56.735 47.785 57.850 ;
		LAYER VIA3 ;
		RECT 47.605 56.405 47.785 56.425 ;
		LAYER M2 ;
		RECT 47.605 55.410 47.785 55.765 ;
		LAYER M3 ;
		RECT 47.605 54.745 47.785 54.765 ;
		LAYER M2 ;
		RECT 47.605 54.415 47.785 54.435 ;
		LAYER M3 ;
		RECT 47.605 54.415 47.785 54.435 ;
		LAYER M1 ;
		RECT 47.605 54.395 47.785 54.455 ;
		LAYER VIA3 ;
		RECT 47.605 54.415 47.785 54.435 ;
		LAYER VIA3 ;
		RECT 47.605 54.745 47.785 54.765 ;
		LAYER M2 ;
		RECT 47.605 50.770 47.785 51.125 ;
		LAYER VIA3 ;
		RECT 47.605 50.770 47.785 51.125 ;
		LAYER M1 ;
		RECT 47.605 53.735 47.785 53.795 ;
		LAYER M2 ;
		RECT 47.605 54.085 47.785 54.105 ;
		LAYER M3 ;
		RECT 47.605 54.085 47.785 54.105 ;
		LAYER VIA3 ;
		RECT 47.605 54.085 47.785 54.105 ;
		LAYER M1 ;
		RECT 47.605 54.065 47.785 54.125 ;
		LAYER M2 ;
		RECT 47.605 48.450 47.785 48.470 ;
		LAYER M1 ;
		RECT 47.605 49.425 47.785 49.485 ;
		LAYER VIA3 ;
		RECT 47.605 49.445 47.785 49.465 ;
		LAYER M1 ;
		RECT 47.605 49.755 47.785 49.815 ;
		LAYER M2 ;
		RECT 47.605 50.105 47.785 50.125 ;
		LAYER M3 ;
		RECT 47.605 50.105 47.785 50.125 ;
		LAYER VIA3 ;
		RECT 47.605 50.105 47.785 50.125 ;
		LAYER M1 ;
		RECT 47.605 48.430 47.785 48.490 ;
		LAYER M1 ;
		RECT 47.605 50.085 47.785 50.145 ;
		LAYER M2 ;
		RECT 47.605 50.435 47.785 50.460 ;
		LAYER M2 ;
		RECT 47.605 46.800 47.785 46.820 ;
		LAYER M1 ;
		RECT 47.605 47.440 47.785 47.500 ;
		LAYER M3 ;
		RECT 47.605 47.460 47.785 47.480 ;
		LAYER M1 ;
		RECT 47.605 50.415 47.785 50.480 ;
		LAYER VIA3 ;
		RECT 47.605 50.435 47.785 50.460 ;
		LAYER M2 ;
		RECT 47.605 49.445 47.785 49.465 ;
		LAYER M3 ;
		RECT 47.605 49.445 47.785 49.465 ;
		LAYER M3 ;
		RECT 47.605 50.435 47.785 50.460 ;
		LAYER M2 ;
		RECT 47.605 49.775 47.785 49.795 ;
		LAYER M3 ;
		RECT 47.605 49.775 47.785 49.795 ;
		LAYER VIA3 ;
		RECT 47.605 49.775 47.785 49.795 ;
		LAYER M3 ;
		RECT 47.605 53.755 47.785 53.775 ;
		LAYER M2 ;
		RECT 47.605 53.090 47.785 53.445 ;
		LAYER M3 ;
		RECT 47.605 53.090 47.785 53.445 ;
		LAYER M1 ;
		RECT 47.605 53.070 47.785 53.465 ;
		LAYER VIA3 ;
		RECT 47.605 53.090 47.785 53.445 ;
		LAYER M2 ;
		RECT 47.605 51.765 47.785 51.785 ;
		LAYER M3 ;
		RECT 47.605 51.765 47.785 51.785 ;
		LAYER VIA3 ;
		RECT 47.605 51.765 47.785 51.785 ;
		LAYER M1 ;
		RECT 47.605 51.745 47.785 51.805 ;
		LAYER M1 ;
		RECT 47.605 52.735 47.785 52.800 ;
		LAYER M3 ;
		RECT 47.605 52.425 47.785 52.445 ;
		LAYER M1 ;
		RECT 47.605 52.405 47.785 52.465 ;
		LAYER M1 ;
		RECT 47.605 50.750 47.785 51.145 ;
		LAYER VIA3 ;
		RECT 47.605 51.435 47.785 51.455 ;
		LAYER M2 ;
		RECT 47.605 51.435 47.785 51.455 ;
		LAYER M1 ;
		RECT 47.605 51.415 47.785 51.475 ;
		LAYER M3 ;
		RECT 47.605 51.435 47.785 51.455 ;
		LAYER M3 ;
		RECT 47.605 50.770 47.785 51.125 ;
		LAYER VIA3 ;
		RECT 47.605 53.755 47.785 53.775 ;
		LAYER M2 ;
		RECT 47.605 52.755 47.785 52.780 ;
		LAYER M3 ;
		RECT 47.605 52.755 47.785 52.780 ;
		LAYER VIA3 ;
		RECT 47.605 52.755 47.785 52.780 ;
		LAYER M1 ;
		RECT 47.605 52.075 47.785 52.135 ;
		LAYER VIA3 ;
		RECT 47.605 52.095 47.785 52.115 ;
		LAYER M3 ;
		RECT 47.605 52.095 47.785 52.115 ;
		LAYER VIA3 ;
		RECT 47.605 52.425 47.785 52.445 ;
		LAYER M2 ;
		RECT 47.605 52.095 47.785 52.115 ;
		LAYER M2 ;
		RECT 47.605 52.425 47.785 52.445 ;
		LAYER M1 ;
		RECT 47.605 46.780 47.785 46.840 ;
		LAYER M2 ;
		RECT 47.605 47.460 47.785 47.480 ;
		LAYER VIA3 ;
		RECT 47.605 47.460 47.785 47.480 ;
		LAYER VIA3 ;
		RECT 47.605 46.800 47.785 46.820 ;
		LAYER M3 ;
		RECT 47.605 46.800 47.785 46.820 ;
		LAYER M2 ;
		RECT 47.605 47.130 47.785 47.150 ;
		LAYER M3 ;
		RECT 47.605 47.130 47.785 47.150 ;
		LAYER VIA3 ;
		RECT 47.605 47.130 47.785 47.150 ;
		LAYER M1 ;
		RECT 47.605 47.110 47.785 47.170 ;
		LAYER M2 ;
		RECT 47.605 47.790 47.785 47.810 ;
		LAYER M3 ;
		RECT 47.605 47.790 47.785 47.810 ;
		LAYER VIA3 ;
		RECT 47.605 47.790 47.785 47.810 ;
		LAYER M1 ;
		RECT 47.605 47.770 47.785 47.830 ;
		LAYER M2 ;
		RECT 47.605 46.470 47.785 46.490 ;
		LAYER M3 ;
		RECT 47.605 48.120 47.785 48.140 ;
		LAYER VIA3 ;
		RECT 47.605 48.120 47.785 48.140 ;
		LAYER M2 ;
		RECT 47.605 48.120 47.785 48.140 ;
		LAYER M3 ;
		RECT 47.605 46.470 47.785 46.490 ;
		LAYER VIA3 ;
		RECT 47.605 46.470 47.785 46.490 ;
		LAYER M1 ;
		RECT 47.605 48.100 47.785 48.160 ;
		LAYER M2 ;
		RECT 47.605 53.755 47.785 53.775 ;
		LAYER VIA3 ;
		RECT 47.605 12.675 47.785 12.695 ;
		LAYER M2 ;
		RECT 47.605 12.675 47.785 12.695 ;
		LAYER M3 ;
		RECT 47.605 12.675 47.785 12.695 ;
		LAYER M2 ;
		RECT 47.605 10.695 47.785 10.715 ;
		LAYER M2 ;
		RECT 47.605 10.365 47.785 10.385 ;
		LAYER M3 ;
		RECT 47.605 10.365 47.785 10.385 ;
		LAYER VIA3 ;
		RECT 47.605 10.365 47.785 10.385 ;
		LAYER M2 ;
		RECT 47.605 8.055 47.785 8.075 ;
		LAYER VIA3 ;
		RECT 47.605 9.375 47.785 9.395 ;
		LAYER M2 ;
		RECT 47.605 9.375 47.785 9.395 ;
		LAYER M2 ;
		RECT 47.605 9.705 47.785 10.055 ;
		LAYER M3 ;
		RECT 47.605 8.055 47.785 8.075 ;
		LAYER M1 ;
		RECT 47.605 9.685 47.785 10.075 ;
		LAYER M3 ;
		RECT 47.605 9.705 47.785 10.055 ;
		LAYER M1 ;
		RECT 47.605 10.345 47.785 10.405 ;
		LAYER M3 ;
		RECT 47.605 11.685 47.785 11.705 ;
		LAYER M3 ;
		RECT 47.605 12.015 47.785 12.035 ;
		LAYER VIA3 ;
		RECT 47.605 12.015 47.785 12.035 ;
		LAYER VIA3 ;
		RECT 47.605 11.685 47.785 11.705 ;
		LAYER M2 ;
		RECT 47.605 11.685 47.785 11.705 ;
		LAYER M1 ;
		RECT 47.605 11.995 47.785 12.055 ;
		LAYER M3 ;
		RECT 47.605 12.345 47.785 12.365 ;
		LAYER VIA3 ;
		RECT 47.605 12.345 47.785 12.365 ;
		LAYER M1 ;
		RECT 47.605 12.325 47.785 12.385 ;
		LAYER M1 ;
		RECT 47.605 40.840 47.785 40.900 ;
		LAYER M1 ;
		RECT 47.605 40.510 47.785 40.570 ;
		LAYER M1 ;
		RECT 47.605 46.450 47.785 46.510 ;
		LAYER M1 ;
		RECT 47.605 37.565 47.785 37.630 ;
		LAYER M2 ;
		RECT 47.605 36.600 47.785 36.620 ;
		LAYER M3 ;
		RECT 47.605 36.600 47.785 36.620 ;
		LAYER M1 ;
		RECT 47.605 36.580 47.785 36.640 ;
		LAYER M1 ;
		RECT 47.605 37.240 47.785 37.295 ;
		LAYER M1 ;
		RECT 47.605 37.900 47.785 37.960 ;
		LAYER M2 ;
		RECT 47.605 37.920 47.785 37.940 ;
		LAYER M1 ;
		RECT 47.605 34.930 47.785 36.310 ;
		LAYER M1 ;
		RECT 47.605 32.985 47.785 34.000 ;
		LAYER M2 ;
		RECT 47.605 33.005 47.785 33.980 ;
		LAYER M2 ;
		RECT 47.605 32.675 47.785 32.695 ;
		LAYER M1 ;
		RECT 47.605 32.655 47.785 32.715 ;
		LAYER M3 ;
		RECT 47.605 11.355 47.785 11.375 ;
		LAYER VIA3 ;
		RECT 47.605 10.695 47.785 10.715 ;
		LAYER M1 ;
		RECT 47.605 10.675 47.785 10.735 ;
		LAYER M2 ;
		RECT 47.605 11.355 47.785 11.375 ;
		LAYER M2 ;
		RECT 47.605 11.025 47.785 11.045 ;
		LAYER M3 ;
		RECT 47.605 11.025 47.785 11.045 ;
		LAYER VIA3 ;
		RECT 47.605 11.025 47.785 11.045 ;
		LAYER M1 ;
		RECT 47.605 11.005 47.785 11.065 ;
		LAYER M1 ;
		RECT 47.605 11.335 47.785 11.395 ;
		LAYER VIA3 ;
		RECT 47.605 11.355 47.785 11.375 ;
		LAYER M3 ;
		RECT 47.605 10.695 47.785 10.715 ;
		LAYER M3 ;
		RECT 47.605 4.410 47.785 4.765 ;
		LAYER VIA3 ;
		RECT 47.605 4.410 47.785 4.765 ;
		LAYER M1 ;
		RECT 47.605 5.385 47.785 5.445 ;
		LAYER M2 ;
		RECT 47.605 5.405 47.785 5.425 ;
		LAYER M3 ;
		RECT 47.605 5.405 47.785 5.425 ;
		LAYER M2 ;
		RECT 47.605 5.735 47.785 5.755 ;
		LAYER M3 ;
		RECT 47.605 5.735 47.785 5.755 ;
		LAYER VIA3 ;
		RECT 47.605 5.735 47.785 5.755 ;
		LAYER VIA3 ;
		RECT 47.605 5.405 47.785 5.425 ;
		LAYER M2 ;
		RECT 47.605 6.065 47.785 6.085 ;
		LAYER M3 ;
		RECT 47.605 6.065 47.785 6.085 ;
		LAYER M1 ;
		RECT 47.605 5.715 47.785 5.775 ;
		LAYER M1 ;
		RECT 47.605 6.045 47.785 6.105 ;
		LAYER VIA3 ;
		RECT 47.605 6.065 47.785 6.085 ;
		LAYER M1 ;
		RECT 47.605 7.375 47.785 7.435 ;
		LAYER VIA3 ;
		RECT 47.605 6.730 47.785 7.085 ;
		LAYER M1 ;
		RECT 47.605 6.710 47.785 7.105 ;
		LAYER VIA3 ;
		RECT 47.605 6.395 47.785 6.420 ;
		LAYER VIA3 ;
		RECT 47.605 7.395 47.785 7.415 ;
		LAYER M2 ;
		RECT 47.605 7.395 47.785 7.415 ;
		LAYER M3 ;
		RECT 47.605 7.395 47.785 7.415 ;
		LAYER M1 ;
		RECT 47.605 6.375 47.785 6.440 ;
		LAYER M2 ;
		RECT 47.605 5.075 47.785 5.095 ;
		LAYER M3 ;
		RECT 47.605 5.075 47.785 5.095 ;
		LAYER VIA3 ;
		RECT 47.605 5.075 47.785 5.095 ;
		LAYER M1 ;
		RECT 47.605 5.055 47.785 5.115 ;
		LAYER M2 ;
		RECT 47.605 6.730 47.785 7.085 ;
		LAYER M1 ;
		RECT 47.605 7.705 47.785 7.765 ;
		LAYER VIA3 ;
		RECT 47.605 7.725 47.785 7.745 ;
		LAYER M2 ;
		RECT 47.605 9.045 47.785 9.065 ;
		LAYER M3 ;
		RECT 47.605 9.045 47.785 9.065 ;
		LAYER VIA3 ;
		RECT 47.605 9.045 47.785 9.065 ;
		LAYER VIA3 ;
		RECT 47.605 8.715 47.785 8.735 ;
		LAYER M2 ;
		RECT 47.605 8.715 47.785 8.735 ;
		LAYER M3 ;
		RECT 47.605 8.715 47.785 8.735 ;
		LAYER M3 ;
		RECT 47.605 6.730 47.785 7.085 ;
		LAYER M1 ;
		RECT 47.605 9.025 47.785 9.085 ;
		LAYER M3 ;
		RECT 47.605 9.375 47.785 9.395 ;
		LAYER M1 ;
		RECT 47.605 9.355 47.785 9.415 ;
		LAYER M1 ;
		RECT 47.605 8.035 47.785 8.095 ;
		LAYER M2 ;
		RECT 47.605 6.395 47.785 6.420 ;
		LAYER M3 ;
		RECT 47.605 6.395 47.785 6.420 ;
		LAYER VIA3 ;
		RECT 47.605 9.705 47.785 10.055 ;
		LAYER VIA3 ;
		RECT 47.605 8.385 47.785 8.405 ;
		LAYER M1 ;
		RECT 47.605 8.365 47.785 8.425 ;
		LAYER VIA3 ;
		RECT 47.605 8.055 47.785 8.075 ;
		LAYER M1 ;
		RECT 47.605 8.695 47.785 8.755 ;
		LAYER M2 ;
		RECT 47.605 56.735 47.785 57.850 ;
		LAYER M1 ;
		RECT 47.605 55.055 47.785 55.120 ;
		LAYER VIA3 ;
		RECT 47.605 55.075 47.785 55.100 ;
		LAYER M2 ;
		RECT 47.605 56.405 47.785 56.425 ;
		LAYER M3 ;
		RECT 47.605 55.075 47.785 55.100 ;
		LAYER M1 ;
		RECT 47.605 55.390 47.785 55.785 ;
		LAYER M3 ;
		RECT 47.605 55.410 47.785 55.765 ;
		LAYER VIA3 ;
		RECT 47.605 55.410 47.785 55.765 ;
		LAYER M2 ;
		RECT 47.605 55.075 47.785 55.100 ;
		LAYER M1 ;
		RECT 47.605 56.385 47.785 56.445 ;
		LAYER M2 ;
		RECT 47.605 56.075 47.785 56.095 ;
		LAYER M3 ;
		RECT 47.605 56.075 47.785 56.095 ;
		LAYER M1 ;
		RECT 47.605 56.055 47.785 56.115 ;
		LAYER VIA3 ;
		RECT 47.605 56.075 47.785 56.095 ;
		LAYER M1 ;
		RECT 47.605 17.530 47.785 17.610 ;
		LAYER M2 ;
		RECT 47.605 16.890 47.785 16.910 ;
		LAYER M2 ;
		RECT 47.605 16.560 47.785 16.580 ;
		LAYER M2 ;
		RECT 47.605 15.900 47.785 15.920 ;
		LAYER M2 ;
		RECT 47.605 16.230 47.785 16.250 ;
		LAYER M3 ;
		RECT 47.605 44.490 47.785 44.510 ;
		LAYER VIA3 ;
		RECT 47.605 44.490 47.785 44.510 ;
		LAYER M1 ;
		RECT 47.605 38.230 47.785 38.290 ;
		LAYER M1 ;
		RECT 47.605 44.470 47.785 44.530 ;
		LAYER M2 ;
		RECT 47.605 44.490 47.785 44.510 ;
		LAYER M1 ;
		RECT 47.605 43.480 47.785 43.870 ;
		LAYER M2 ;
		RECT 47.605 44.160 47.785 44.180 ;
		LAYER M3 ;
		RECT 47.605 44.160 47.785 44.180 ;
		LAYER M1 ;
		RECT 47.605 44.140 47.785 44.200 ;
		LAYER VIA3 ;
		RECT 47.605 44.160 47.785 44.180 ;
		LAYER M1 ;
		RECT 47.605 22.555 47.785 23.075 ;
		LAYER M1 ;
		RECT 47.605 23.345 47.785 23.405 ;
		LAYER M2 ;
		RECT 47.605 23.365 47.785 23.385 ;
		LAYER M2 ;
		RECT 47.605 22.575 47.785 23.055 ;
		LAYER M3 ;
		RECT 47.605 22.575 47.785 23.055 ;
		LAYER VIA3 ;
		RECT 47.605 22.575 47.785 23.055 ;
		LAYER M2 ;
		RECT 47.605 17.900 47.785 17.920 ;
		LAYER VIA3 ;
		RECT 47.605 18.230 47.785 18.295 ;
		LAYER M2 ;
		RECT 47.605 18.605 47.785 18.625 ;
		LAYER M1 ;
		RECT 47.605 18.585 47.785 18.645 ;
		LAYER VIA3 ;
		RECT 47.605 18.935 47.785 18.955 ;
		LAYER M1 ;
		RECT 47.605 15.220 47.785 15.280 ;
		LAYER M1 ;
		RECT 47.605 15.550 47.785 15.610 ;
		LAYER M2 ;
		RECT 47.605 13.665 47.785 13.685 ;
		LAYER M3 ;
		RECT 47.605 13.665 47.785 13.685 ;
		LAYER M1 ;
		RECT 47.605 13.645 47.785 13.705 ;
		LAYER M3 ;
		RECT 47.605 13.995 47.785 14.930 ;
		LAYER VIA3 ;
		RECT 47.605 13.665 47.785 13.685 ;
		LAYER VIA3 ;
		RECT 47.605 13.995 47.785 14.930 ;
		LAYER M3 ;
		RECT 47.605 15.240 47.785 15.260 ;
		LAYER VIA3 ;
		RECT 47.605 15.240 47.785 15.260 ;
		LAYER M2 ;
		RECT 47.605 15.240 47.785 15.260 ;
		LAYER M2 ;
		RECT 47.605 13.995 47.785 14.930 ;
		LAYER M2 ;
		RECT 47.605 40.860 47.785 40.880 ;
		LAYER M3 ;
		RECT 47.605 40.860 47.785 40.880 ;
		LAYER M3 ;
		RECT 47.605 41.190 47.785 41.210 ;
		LAYER M2 ;
		RECT 47.605 41.190 47.785 41.210 ;
		LAYER VIA3 ;
		RECT 47.605 41.190 47.785 41.210 ;
		LAYER VIA3 ;
		RECT 47.605 40.860 47.785 40.880 ;
		LAYER M1 ;
		RECT 47.605 42.490 47.785 42.550 ;
		LAYER M1 ;
		RECT 47.605 41.170 47.785 41.230 ;
		LAYER M1 ;
		RECT 47.605 41.500 47.785 41.560 ;
		LAYER M3 ;
		RECT 47.605 43.170 47.785 43.190 ;
		LAYER M2 ;
		RECT 47.605 43.500 47.785 43.850 ;
		LAYER M3 ;
		RECT 47.605 43.500 47.785 43.850 ;
		LAYER VIA3 ;
		RECT 47.605 43.500 47.785 43.850 ;
		LAYER M1 ;
		RECT 47.605 43.150 47.785 43.210 ;
		LAYER M3 ;
		RECT 47.605 41.850 47.785 42.200 ;
		LAYER VIA3 ;
		RECT 47.605 41.850 47.785 42.200 ;
		LAYER M2 ;
		RECT 47.605 41.850 47.785 42.200 ;
		LAYER M1 ;
		RECT 47.605 41.830 47.785 42.220 ;
		LAYER M2 ;
		RECT 47.605 41.520 47.785 41.540 ;
		LAYER VIA3 ;
		RECT 47.605 41.520 47.785 41.540 ;
		LAYER M3 ;
		RECT 47.605 41.520 47.785 41.540 ;
		LAYER M1 ;
		RECT 47.605 42.820 47.785 42.880 ;
		LAYER M2 ;
		RECT 47.605 42.510 47.785 42.530 ;
		LAYER M3 ;
		RECT 47.605 42.510 47.785 42.530 ;
		LAYER VIA3 ;
		RECT 47.605 42.510 47.785 42.530 ;
		LAYER M2 ;
		RECT 47.605 43.170 47.785 43.190 ;
		LAYER M2 ;
		RECT 47.605 42.840 47.785 42.860 ;
		LAYER M3 ;
		RECT 47.605 42.840 47.785 42.860 ;
		LAYER VIA3 ;
		RECT 47.605 42.840 47.785 42.860 ;
		LAYER VIA3 ;
		RECT 47.605 43.170 47.785 43.190 ;
		LAYER M2 ;
		RECT 47.605 23.695 47.785 23.745 ;
		LAYER M1 ;
		RECT 47.605 23.675 47.785 23.765 ;
		LAYER M2 ;
		RECT 47.605 24.055 47.785 24.075 ;
		LAYER M3 ;
		RECT 47.605 24.055 47.785 24.075 ;
		LAYER M3 ;
		RECT 47.605 23.695 47.785 23.745 ;
		LAYER VIA3 ;
		RECT 47.605 23.695 47.785 23.745 ;
		LAYER M1 ;
		RECT 47.605 12.985 47.785 13.045 ;
		LAYER M1 ;
		RECT 47.605 13.975 47.785 14.950 ;
		LAYER M2 ;
		RECT 47.605 13.005 47.785 13.025 ;
		LAYER M3 ;
		RECT 47.605 13.005 47.785 13.025 ;
		LAYER VIA3 ;
		RECT 47.605 13.005 47.785 13.025 ;
		LAYER M1 ;
		RECT 47.605 13.315 47.785 13.375 ;
		LAYER M2 ;
		RECT 47.605 13.335 47.785 13.355 ;
		LAYER M3 ;
		RECT 47.605 13.335 47.785 13.355 ;
		LAYER VIA3 ;
		RECT 47.605 13.335 47.785 13.355 ;
		LAYER M1 ;
		RECT 47.605 17.880 47.785 17.940 ;
		LAYER M2 ;
		RECT 47.605 18.935 47.785 18.955 ;
		LAYER M1 ;
		RECT 47.605 19.245 47.785 21.955 ;
		LAYER M1 ;
		RECT 47.605 38.560 47.785 38.620 ;
		LAYER M1 ;
		RECT 47.605 24.365 47.785 29.505 ;
		LAYER M2 ;
		RECT 47.605 24.385 47.785 29.485 ;
		LAYER M1 ;
		RECT 47.605 24.035 47.785 24.095 ;
		LAYER M3 ;
		RECT 47.605 37.920 47.785 37.940 ;
		LAYER VIA3 ;
		RECT 47.605 37.920 47.785 37.940 ;
		LAYER M1 ;
		RECT 47.605 36.910 47.785 36.970 ;
		LAYER VIA3 ;
		RECT 47.605 36.600 47.785 36.620 ;
		LAYER M2 ;
		RECT 47.605 34.950 47.785 36.290 ;
		LAYER M3 ;
		RECT 47.605 34.950 47.785 36.290 ;
		LAYER M2 ;
		RECT 47.605 29.795 47.785 29.815 ;
		LAYER M3 ;
		RECT 47.605 29.795 47.785 29.815 ;
		LAYER M1 ;
		RECT 47.605 30.105 47.785 31.725 ;
		LAYER VIA3 ;
		RECT 47.605 29.795 47.785 29.815 ;
		LAYER M1 ;
		RECT 47.605 29.775 47.785 29.835 ;
		LAYER VIA3 ;
		RECT 47.605 24.385 47.785 29.485 ;
		LAYER M3 ;
		RECT 47.605 24.385 47.785 29.485 ;
		LAYER M1 ;
		RECT 47.605 40.180 47.785 40.240 ;
		LAYER M3 ;
		RECT 47.605 40.200 47.785 40.220 ;
		LAYER M1 ;
		RECT 47.605 39.220 47.785 39.910 ;
		LAYER M2 ;
		RECT 47.605 38.580 47.785 38.600 ;
		LAYER M2 ;
		RECT 47.605 34.620 47.785 34.640 ;
		LAYER M1 ;
		RECT 47.605 34.270 47.785 34.330 ;
		LAYER M3 ;
		RECT 47.605 33.005 47.785 33.980 ;
		LAYER VIA3 ;
		RECT 47.605 33.005 47.785 33.980 ;
		LAYER M3 ;
		RECT 47.605 32.675 47.785 32.695 ;
		LAYER VIA3 ;
		RECT 47.605 32.675 47.785 32.695 ;
		LAYER M1 ;
		RECT 47.605 34.600 47.785 34.660 ;
		LAYER M2 ;
		RECT 47.605 34.290 47.785 34.310 ;
		LAYER VIA3 ;
		RECT 47.605 34.290 47.785 34.310 ;
		LAYER M3 ;
		RECT 47.605 34.290 47.785 34.310 ;
		LAYER M3 ;
		RECT 47.605 32.345 47.785 32.365 ;
		LAYER M3 ;
		RECT 47.605 32.015 47.785 32.035 ;
		LAYER VIA3 ;
		RECT 47.605 32.015 47.785 32.035 ;
		LAYER M2 ;
		RECT 47.605 32.015 47.785 32.035 ;
		LAYER M1 ;
		RECT 47.605 32.325 47.785 32.385 ;
		LAYER M2 ;
		RECT 47.605 32.345 47.785 32.365 ;
		LAYER VIA3 ;
		RECT 47.605 32.345 47.785 32.365 ;
		LAYER M2 ;
		RECT 47.605 30.125 47.785 31.705 ;
		LAYER M1 ;
		RECT 47.605 31.995 47.785 32.055 ;
		LAYER M3 ;
		RECT 47.605 30.125 47.785 31.705 ;
		LAYER VIA3 ;
		RECT 47.605 30.125 47.785 31.705 ;
		LAYER M2 ;
		RECT 47.605 40.530 47.785 40.550 ;
		LAYER M2 ;
		RECT 47.605 40.200 47.785 40.220 ;
		LAYER VIA3 ;
		RECT 47.605 40.200 47.785 40.220 ;
		LAYER VIA3 ;
		RECT 47.605 40.530 47.785 40.550 ;
		LAYER M3 ;
		RECT 47.605 40.530 47.785 40.550 ;
		LAYER M3 ;
		RECT 47.605 34.620 47.785 34.640 ;
		LAYER VIA3 ;
		RECT 47.605 34.620 47.785 34.640 ;
		LAYER VIA3 ;
		RECT 47.605 34.950 47.785 36.290 ;
		LAYER VIA3 ;
		RECT 47.605 39.240 47.785 39.890 ;
		LAYER M2 ;
		RECT 47.605 39.240 47.785 39.890 ;
		LAYER M3 ;
		RECT 47.605 39.240 47.785 39.890 ;
		LAYER M1 ;
		RECT 47.605 38.890 47.785 38.950 ;
		LAYER M2 ;
		RECT 47.605 22.245 47.785 22.265 ;
		LAYER M1 ;
		RECT 47.605 22.225 47.785 22.285 ;
		LAYER M2 ;
		RECT 47.605 19.265 47.785 21.935 ;
		LAYER M3 ;
		RECT 47.605 19.265 47.785 21.935 ;
		LAYER M2 ;
		RECT 47.605 17.550 47.785 17.590 ;
		LAYER M3 ;
		RECT 47.605 17.900 47.785 17.920 ;
		LAYER M2 ;
		RECT 47.605 18.230 47.785 18.295 ;
		LAYER M3 ;
		RECT 47.605 18.230 47.785 18.295 ;
		LAYER M1 ;
		RECT 47.605 17.200 47.785 17.260 ;
		LAYER M3 ;
		RECT 47.605 17.220 47.785 17.240 ;
		LAYER M1 ;
		RECT 47.605 16.540 47.785 16.600 ;
		LAYER M2 ;
		RECT 47.605 17.220 47.785 17.240 ;
		LAYER VIA3 ;
		RECT 47.605 17.220 47.785 17.240 ;
		LAYER VIA3 ;
		RECT 47.605 17.900 47.785 17.920 ;
		LAYER M1 ;
		RECT 47.605 16.210 47.785 16.270 ;
		LAYER VIA3 ;
		RECT 47.605 16.230 47.785 16.250 ;
		LAYER M3 ;
		RECT 47.605 16.890 47.785 16.910 ;
		LAYER VIA3 ;
		RECT 47.605 16.890 47.785 16.910 ;
		LAYER M1 ;
		RECT 47.605 16.870 47.785 16.930 ;
		LAYER M3 ;
		RECT 47.605 16.560 47.785 16.580 ;
		LAYER VIA3 ;
		RECT 47.605 16.560 47.785 16.580 ;
		LAYER M3 ;
		RECT 47.605 17.550 47.785 17.590 ;
		LAYER VIA3 ;
		RECT 47.605 17.550 47.785 17.590 ;
		LAYER VIA3 ;
		RECT 47.605 18.605 47.785 18.625 ;
		LAYER M1 ;
		RECT 47.605 18.210 47.785 18.315 ;
		LAYER M3 ;
		RECT 47.605 22.245 47.785 22.265 ;
		LAYER VIA3 ;
		RECT 47.605 22.245 47.785 22.265 ;
		LAYER VIA3 ;
		RECT 47.605 19.265 47.785 21.935 ;
		LAYER VIA3 ;
		RECT 47.605 24.055 47.785 24.075 ;
		LAYER M1 ;
		RECT 47.605 18.915 47.785 18.975 ;
		LAYER M3 ;
		RECT 47.605 18.935 47.785 18.955 ;
		LAYER M3 ;
		RECT 47.605 23.365 47.785 23.385 ;
		LAYER VIA3 ;
		RECT 47.605 23.365 47.785 23.385 ;
		LAYER M3 ;
		RECT 47.605 18.605 47.785 18.625 ;
		LAYER M2 ;
		RECT 47.605 15.570 47.785 15.590 ;
		LAYER M3 ;
		RECT 47.605 15.570 47.785 15.590 ;
		LAYER VIA3 ;
		RECT 47.605 15.570 47.785 15.590 ;
		LAYER M3 ;
		RECT 47.605 15.900 47.785 15.920 ;
		LAYER VIA3 ;
		RECT 47.605 15.900 47.785 15.920 ;
		LAYER M1 ;
		RECT 47.605 15.880 47.785 15.940 ;
		LAYER M3 ;
		RECT 47.605 16.230 47.785 16.250 ;
		LAYER M2 ;
		RECT 47.605 38.250 47.785 38.270 ;
		LAYER M3 ;
		RECT 47.605 38.250 47.785 38.270 ;
		LAYER VIA3 ;
		RECT 47.605 38.250 47.785 38.270 ;
		LAYER M3 ;
		RECT 47.605 38.580 47.785 38.600 ;
		LAYER M2 ;
		RECT 47.605 38.910 47.785 38.930 ;
		LAYER M3 ;
		RECT 47.605 38.910 47.785 38.930 ;
		LAYER VIA3 ;
		RECT 47.605 38.910 47.785 38.930 ;
		LAYER M2 ;
		RECT 47.605 37.585 47.785 37.610 ;
		LAYER M3 ;
		RECT 47.605 37.585 47.785 37.610 ;
		LAYER VIA3 ;
		RECT 47.605 37.585 47.785 37.610 ;
		LAYER VIA3 ;
		RECT 47.605 38.580 47.785 38.600 ;
		LAYER VIA3 ;
		RECT 47.605 36.930 47.785 36.950 ;
		LAYER M2 ;
		RECT 47.605 36.930 47.785 36.950 ;
		LAYER M3 ;
		RECT 47.605 36.930 47.785 36.950 ;
		LAYER M2 ;
		RECT 47.605 37.260 47.785 37.275 ;
		LAYER VIA3 ;
		RECT 47.605 37.260 47.785 37.275 ;
		LAYER M3 ;
		RECT 47.605 37.260 47.785 37.275 ;
		LAYER M4 ;
		RECT 24.150 29.050 47.395 29.480 ;
		LAYER M4 ;
		RECT 21.525 23.090 47.395 23.850 ;
		LAYER M4 ;
		RECT 21.525 20.290 47.395 22.310 ;
		LAYER M4 ;
		RECT 0.000 24.400 47.395 24.905 ;
		LAYER M4 ;
		RECT 0.000 20.290 21.525 23.850 ;
		LAYER M4 ;
		RECT 0.000 45.765 47.395 46.845 ;
		LAYER M4 ;
		RECT 0.000 48.085 47.395 49.165 ;
		LAYER M3 ;
		RECT 0.000 0.000 47.605 57.850 ;
		LAYER M4 ;
		RECT 0.000 43.445 47.395 44.525 ;
		LAYER M4 ;
		RECT 0.000 41.125 47.395 42.205 ;
		LAYER M4 ;
		RECT 0.000 38.805 47.395 39.885 ;
		LAYER M2 ;
		RECT 0.000 0.000 47.605 57.850 ;
		LAYER M1 ;
		RECT 47.605 12.655 47.785 12.715 ;
		LAYER M1 ;
		RECT 47.605 11.665 47.785 11.725 ;
		LAYER M2 ;
		RECT 47.605 12.345 47.785 12.365 ;
		LAYER M2 ;
		RECT 47.605 12.015 47.785 12.035 ;
		LAYER M1 ;
		RECT 47.605 0.000 47.785 1.135 ;
		LAYER M3 ;
		RECT 47.605 0.000 47.785 1.115 ;
		LAYER VIA3 ;
		RECT 47.605 0.000 47.785 1.115 ;
		LAYER VIA3 ;
		RECT 47.605 2.090 47.785 2.445 ;
		LAYER M3 ;
		RECT 47.605 2.090 47.785 2.445 ;
		LAYER M1 ;
		RECT 47.605 2.070 47.785 2.465 ;
		LAYER M1 ;
		RECT 47.605 1.735 47.785 1.800 ;
		LAYER M2 ;
		RECT 47.605 2.090 47.785 2.445 ;
		LAYER M2 ;
		RECT 47.605 0.000 47.785 1.115 ;
		LAYER M2 ;
		RECT 47.605 1.755 47.785 1.780 ;
		LAYER VIA3 ;
		RECT 47.605 1.755 47.785 1.780 ;
		LAYER M3 ;
		RECT 47.605 1.755 47.785 1.780 ;
		LAYER M3 ;
		RECT 47.605 1.425 47.785 1.445 ;
		LAYER M2 ;
		RECT 47.605 1.425 47.785 1.445 ;
		LAYER VIA3 ;
		RECT 47.605 1.425 47.785 1.445 ;
		LAYER M1 ;
		RECT 47.605 1.405 47.785 1.465 ;
		LAYER M4 ;
		RECT 0.000 55.045 47.395 56.125 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 47.785 57.850 ;
		LAYER M1 ;
		RECT 0.000 0.000 47.605 57.850 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 47.785 57.850 ;
		LAYER M1 ;
		RECT 47.605 2.735 47.785 2.795 ;
		LAYER M2 ;
		RECT 47.605 2.755 47.785 2.775 ;
		LAYER M1 ;
		RECT 47.605 4.390 47.785 4.785 ;
		LAYER M3 ;
		RECT 47.605 2.755 47.785 2.775 ;
		LAYER VIA3 ;
		RECT 47.605 2.755 47.785 2.775 ;
		LAYER M1 ;
		RECT 47.605 3.725 47.785 3.785 ;
		LAYER VIA3 ;
		RECT 47.605 4.075 47.785 4.100 ;
		LAYER M2 ;
		RECT 47.605 4.075 47.785 4.100 ;
		LAYER M3 ;
		RECT 47.605 4.075 47.785 4.100 ;
		LAYER VIA3 ;
		RECT 47.605 3.745 47.785 3.765 ;
		LAYER M2 ;
		RECT 47.605 7.725 47.785 7.745 ;
		LAYER M3 ;
		RECT 47.605 7.725 47.785 7.745 ;
		LAYER M2 ;
		RECT 47.605 8.385 47.785 8.405 ;
		LAYER M3 ;
		RECT 47.605 8.385 47.785 8.405 ;
		LAYER M1 ;
		RECT 47.605 3.065 47.785 3.125 ;
		LAYER M2 ;
		RECT 47.605 3.085 47.785 3.105 ;
		LAYER M3 ;
		RECT 47.605 3.085 47.785 3.105 ;
		LAYER M2 ;
		RECT 47.605 4.410 47.785 4.765 ;
		LAYER VIA3 ;
		RECT 47.605 3.085 47.785 3.105 ;
		LAYER M3 ;
		RECT 47.605 3.415 47.785 3.435 ;
		LAYER VIA3 ;
		RECT 47.605 3.415 47.785 3.435 ;
		LAYER M1 ;
		RECT 47.605 3.395 47.785 3.455 ;
		LAYER M2 ;
		RECT 47.605 3.415 47.785 3.435 ;
		LAYER M3 ;
		RECT 47.605 3.745 47.785 3.765 ;
		LAYER M2 ;
		RECT 47.605 3.745 47.785 3.765 ;
		LAYER M1 ;
		RECT 47.605 4.055 47.785 4.120 ;
		LAYER M4 ;
		RECT 0.000 19.425 47.395 19.985 ;
		LAYER M4 ;
		RECT 0.000 15.645 47.395 16.725 ;
		LAYER M4 ;
		RECT 0.000 13.325 47.395 14.405 ;
		LAYER M4 ;
		RECT 24.150 30.930 47.395 31.310 ;
		LAYER M4 ;
		RECT 0.000 29.050 24.150 31.310 ;
		LAYER M4 ;
		RECT 0.000 17.965 47.395 19.045 ;
		LAYER M4 ;
		RECT 0.000 32.680 47.395 34.825 ;
		LAYER M4 ;
		RECT 0.000 11.005 47.395 12.085 ;
		LAYER M4 ;
		RECT 0.000 8.685 47.395 9.765 ;
		LAYER M4 ;
		RECT 0.000 6.365 47.395 7.445 ;
		LAYER M4 ;
		RECT 0.000 35.935 47.395 38.475 ;
		LAYER M4 ;
		RECT 0.000 4.045 47.395 5.125 ;
		LAYER M4 ;
		RECT 0.000 1.725 47.395 2.805 ;
		LAYER M4 ;
		RECT 0.000 52.725 47.395 53.805 ;
		LAYER M4 ;
		RECT 0.000 50.405 47.395 51.485 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 47.605 57.850 ;
	END
	# End of OBS

END TSDN28HPCPUHDB32X16M4MWA

END LIBRARY
