# DESIGN RULE DOCUMENT: T-N28-CL-DR-001 V1.7
# DESIGN RULE DOCUMENT: T-N28-CL-DR-002 V1.5
# P&R TECHNOLOGY FILE VERSION: T-N28-CL-PR-002-E1 V1.5a

#+Note:
#+      1. Please use EDI v14.25-s034 (or later version) for advanced rule modeling support.
#+      2. Antenna ratio defined in OXIDE2 is for OD18.
#+      3. Please use Captable / QRC(recommendation)  to get the accurate RC values.
#+      4. Set the following command in Encounter to get the correct RC values from 
#+         Captable when executing NanoRoute.
#+         setNanoRouteMode -envResistanceFromCapTable true
#+      5. Using TSMC utility for dummy fill is strongly recommended.
#+      6. User can add/remove any preferred viadevice in this tech LEF.
#+Revision Histroy:
#+      1. 20101117 MxLPC rules
#+      2. 20101122 new VIAy.S.3 & My.S.8 rules
#+      3. 20110209 add DFM v01 VMA/HOOK/CAP rule
#+      4. 20110318 refine value in VMA/HOOK/CAP syntax
#+      5. 20110401 Remove VIAx.S.6 & VIAx.S.7
#+      6. 20110401 New viadevice apply VIAx.EN.14 & VIAx.EN.15
#+      7. 20110627 Rectangular VIA for powerplan
#+      8. 20110627 Bridge rule support
#+      9. 20110627 Enhanced Hook rule for M1/M2
#+     10. 20110831 Add 4cut viadevice for wide metal routing
#+     11. 20110921 Update Antenna modeling for top Mu layer
#+     12. 20111108 Enhancement for EFP.VIAx.S.1~6
#+     13. 20111108 New support for Mx.S.37R/VIAx.R.10R/EFP.Mx.EN.1R
#+     14. 20120305 DFM via revision
#+                  *FBD20*,*FBD30*,*PBDB*,*PBDU*,*PBDE*,*FBS25*,*PBSB*,*PBSU*
#+     15. 20120305 RV 2x2 is only allowed in plymide process
#+                  Please refer to v1.2 design rule RV.W.1 
#+                  Set RV default size as 3um x 3um in this TF
#+                  If RV 2x2 is required, please let it unmarked, and let RV 3x3 marked                                    
#+     16. 20130103 Add enhanced Mx.S.8
#+     17. 20130604 Add implant layer VT*
#+     18. 20130807 MINIMUMCUT coding apply LEF58 format in Mx layer for ENCLF-295 elimination
#+     19. 20140516 Update RMS/PEAK EM
#+     20. 20150713 Turn off bridge rules, BR.S1 BR.S2 BR.S3
#+     21. 20150713 New support "LEF58_ENCLOSURE"


VERSION 5.7 ;
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ;

CLEARANCEMEASURE EUCLIDEAN ;
USEMINSPACING OBS OFF ;

UNITS
    CAPACITANCE PICOFARADS 10 ;
    CURRENT MILLIAMPS 10000 ;
    VOLTAGE VOLTS 1000 ;
    FREQUENCY MEGAHERTZ 10 ;
    DATABASE MICRONS 2000 ;
END UNITS

PROPERTYDEFINITIONS
    LIBRARY LEF58_MAXVIASTACK STRING "MAXVIASTACK 4 NOSINGLE RANGE M1 M6 ;" ;
    LAYER LEF58_AREA STRING ;
    LAYER LEF58_ENCLOSURE STRING ;
    LAYER LEF58_SPACING STRING ;
    LAYER LEF58_CUTCLASS STRING ;
    LAYER LEF58_ENCLOSUREEDGE STRING ;
    LAYER LEF58_SPACINGNOTCHLENGTH STRING ;
    LAYER LEF58_SPACINGENDOFNOTCHWIDTH STRING ;
    LAYER LEF58_MINSTEP STRING ;
    LAYER LEF58_SPACINGTABLE STRING ;
    LAYER LEF58_EOLSPACING STRING ;
    #LAYER LEF58_STEPHEIGHT STRING ;
    LAYER LEF58_CORNERFILLSPACING STRING ;
    LAYER LEF58_EOLENCLOSURE STRING ;
    LAYER LEF58_MINIMUMCUT STRING ;
END PROPERTYDEFINITIONS

MANUFACTURINGGRID 0.005000 ;

SITE core
    SIZE 0.135000 BY 0.900000 ; 
    CLASS CORE ;
    SYMMETRY Y ;
END core

SITE bcore
    SIZE 0.135000 BY 1.800000 ; 
    CLASS CORE ;
    SYMMETRY Y ;
END bcore

SITE ccore
    SIZE 0.135000 BY 2.700000 ; 
    CLASS CORE ;
    SYMMETRY Y ;
END ccore

SITE dcore
    SIZE 0.135000 BY 3.600000 ; 
    CLASS CORE ;
    SYMMETRY Y ;
END dcore

SITE gacore
    SIZE 0.540000 BY 0.900000 ; 
    CLASS CORE ;
    SYMMETRY Y ;
END gacore

LAYER PO
    TYPE MASTERSLICE ;
END PO

LAYER CO
    TYPE CUT ;
    PROPERTY LEF58_ENCLOSUREEDGE "ENCLOSUREEDGE ABOVE 0.015 WIDTH 0.08 PARALLEL 0.18 WITHIN 0.06 ;" ;

    ENCLOSURE ABOVE 0 0.02 ;
    ENCLOSURE ABOVE 0.02 0 ;
    ENCLOSURE ABOVE 0 0.03 WIDTH 0.701 ;
    ENCLOSURE ABOVE 0.03 0 WIDTH 0.701 ;
    ENCLOSURE ABOVE 0.015 0.015 ;

END CO

LAYER VTUL_N
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTUL_N
    
LAYER VTUL_P
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTUL_P

LAYER VTL_N
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTL_N

LAYER VTL_P
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTL_P 

LAYER VTH_N
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTH_N

LAYER VTH_P
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTH_P

LAYER VTUH_N
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTUH_N
    
LAYER VTUH_P
    TYPE IMPLANT ;
    WIDTH 0.27 ;
    SPACING 0.27 ;
END VTUH_P

LAYER M1
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.135 0.100 ;
    OFFSET 0.065 0.000 ;
    MINWIDTH 0.050000 ;
    MAXWIDTH 4.500000 ;
    WIDTH 0.050000 ;

    AREA 0.011500 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.050000 MAXEDGES 1 ;
    PROPERTY LEF58_MINSTEP "MINSTEP 0.05 MAXEDGES 1 MINADJACENTLENGTH 0.065 CONVEXCORNER ;" ;
    PROPERTY LEF58_AREA "AREA 0.014000 EXCEPTEDGELENGTH 0.130000 0.200000 EXCEPTMINSIZE 0.050000 0.200000 ;" ;
    PROPERTY LEF58_AREA "AREA 0.038000 EXCEPTEDGELENGTH 0.130000 EXCEPTMINSIZE 0.050000 0.130000 ;" ;

#---RR:RE:EFP.Mx.S.3 hook v01---#
    PROPERTY LEF58_SPACING "
    SPACING 0.07 NOTCHLENGTH 0.155 CONCAVEENDS 0.055 ; " ;

    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.220000  0.470000  0.630000  1.500000
      WIDTH  0.000000  0.050000  0.050000  0.050000  0.050000  0.050000
      WIDTH  0.100000  0.050000  0.060000  0.060000  0.060000  0.060000
      WIDTH  0.180000  0.050000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.470000  0.050000  0.100000  0.130000  0.130000  0.130000
      WIDTH  0.630000  0.050000  0.100000  0.130000  0.150000  0.150000
      WIDTH  1.500000  0.050000  0.100000  0.130000  0.150000  0.500000 ;

#---WMJ---#
    PROPERTY LEF58_SPACINGTABLE "
       SPACINGTABLE JOGTOJOGSPACING 0.3 JOGWIDTH 0.22
       SHORTJOGSPACING 0.06
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.29 LONGJOGSPACING 0.08
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.19 LONGJOGSPACING 0.10
       WIDTH 0.47 PARALLEL 0.5 WITHIN 0.32 LONGJOGSPACING 0.13
       WIDTH 0.63 PARALLEL 0.7 WITHIN 0.34 LONGJOGSPACING 0.15
       WIDTH 1.50 PARALLEL 1.5 WITHIN 0.50 LONGJOGSPACING 0.30 ; " ;

    PROPERTY LEF58_SPACING "
        SPACING 0.060 ENDOFLINE 0.070 WITHIN 0.025 ;
        SPACING 0.070 ENDOFLINE 0.070 WITHIN 0.025 PARALLELEDGE SUBTRACTEOLWIDTH 0.120 WITHIN 0.070 MINLENGTH 0.050 ; " ;

    #MxLPC: Cap Rule 
    PROPERTY LEF58_SPACING "
	SPACING 0.115 ENDOFLINE 0.055 WITHIN 0.000 PARALLELEDGE 0.060 WITHIN 0.120 MINLENGTH 0.150 TWOEDGES SAMEMETAL ; " ;

#    #  BR.S1 BR.S2 BR.S3  #
#    PROPERTY LEF58_SPACING "
#      SPACING 0.236 CONVEXCORNERS EXTENSION 0.16 0.23 ;
#      SPACING 0.080 CONVEXCORNERS EXTENSION 0.23 0.075 SINGLE 0.3 0.08 0.12 SPANLENGTH 0.3 OPPOSITEWIDTH 0.055 OPPOSITEEXTENSION 0.055 0.025 0.1 ;
#      SPACING 0.051 CONVEXCORNERS EXTENSION 0.160 0.115 SAMESIDE 0.09 ; " ;

    PROPERTY LEF58_MINIMUMCUT "
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 WITHIN 0.100000 FROMABOVE ;
    MINIMUMCUT CUTCLASS VSINGLECUT 4 CUTCLASS VDOUBLECUT 2 WIDTH 0.440000 FROMABOVE ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 FROMABOVE LENGTH 0.180000 WITHIN 1.651000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.000000 FROMABOVE LENGTH 1.000000 WITHIN 4.001000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.500000 FROMABOVE LENGTH 5.000000 WITHIN 10.001000 ; " ;

    HEIGHT 0.365 ;
    THICKNESS 0.090000 ;
    FILLACTIVESPACING 0.2 ;
    RESISTANCE RPERSQ 0.407 ;
    CAPACITANCE CPERSQDIST 0.0002 ;
    EDGECAPACITANCE 8.29E-05 ;

    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 17.473521 15.713983 14.571726 14.569677 11.880775 11.005008 10.501241 10.198232 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 70.748390 73.275119 74.116113 37.058681 37.648251 37.774587 37.837755 37.872849 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

END M1

LAYER VIA1
    TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
        CUTCLASS VSINGLECUT WIDTH 0.05 LENGTH 0.05 CUTS 1 ;
        CUTCLASS VDOUBLECUT WIDTH 0.05 LENGTH 0.13 CUTS 2 ;" ;

    #EFP.VIAx.S.1~6
    PROPERTY LEF58_EOLSPACING "
        EOLSPACING 0.08 0.09 CUTCLASS VSINGLECUT TO VDOUBLECUT 0.085 0.09 ENDWIDTH 0.07 PRL -0.04
        ENCLOSURE 0.04 0.00 EXTENSION 0.065 0.12 SPANLENGTH 0.055 ; " ;

    PROPERTY LEF58_SPACINGTABLE "
    	SPACINGTABLE PRL -0.04 MAXXY 
    	CUTCLASS	VSINGLECUT	VDOUBLECUT
    	VSINGLECUT	0.070 0.080	0.075 0.080
    	VDOUBLECUT	0.075 0.080	0.080 0.080 ;" ;

    #Enhanced Mx.S.8
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VSINGLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VDOUBLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;

    

    
    PROPERTY LEF58_ENCLOSUREEDGE "
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ; 
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
	ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1  ;
        ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1 ; " ;
        
 
    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS VSINGLECUT 0 0.03 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.02 0.02 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.01 0.025 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.02 SIDE 0.02 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.03 SIDE 0.01 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.01 SIDE 0.03 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.04 SIDE 0 ;
        " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ;
    DCCURRENTDENSITY	AVERAGE
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ; 

END VIA1

LAYER M2
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.100 0.100 ;
    OFFSET 0.000 0.000 ;
    MINWIDTH 0.050000 ;
    MAXWIDTH 4.500000 ;
    WIDTH 0.050000 ;

    AREA 0.014 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.050000 MAXEDGES 1 ;
    PROPERTY LEF58_MINSTEP "MINSTEP 0.05 MAXEDGES 1 MINADJACENTLENGTH 0.065 CONVEXCORNER ;" ;
    PROPERTY LEF58_AREA "AREA 0.044000 EXCEPTEDGELENGTH 0.130000 EXCEPTMINSIZE 0.050000 0.130000 ;" ;

    #---RR:RE:EFP.Mx.S.3 hook v01---#
    PROPERTY LEF58_SPACING "
    SPACING 0.07 NOTCHLENGTH 0.155 CONCAVEENDS 0.055 ; " ;


    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.220000  0.470000  0.630000  1.500000
      WIDTH  0.000000  0.050000  0.050000  0.050000  0.050000  0.050000
      WIDTH  0.090000  0.050000  0.060000  0.060000  0.060000  0.060000
      WIDTH  0.130000  0.050000  0.080000  0.080000  0.080000  0.080000
      WIDTH  0.160000  0.050000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.470000  0.050000  0.100000  0.130000  0.130000  0.130000
      WIDTH  0.630000  0.050000  0.100000  0.130000  0.150000  0.150000
      WIDTH  1.500000  0.050000  0.100000  0.130000  0.150000  0.500000 ;
    
    PROPERTY LEF58_SPACINGTABLE "
       SPACINGTABLE JOGTOJOGSPACING 0.3 JOGWIDTH 0.22
       SHORTJOGSPACING 0.06
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.29 LONGJOGSPACING 0.08
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.19 LONGJOGSPACING 0.10
       WIDTH 0.47 PARALLEL 0.5 WITHIN 0.32 LONGJOGSPACING 0.13
       WIDTH 0.63 PARALLEL 0.7 WITHIN 0.34 LONGJOGSPACING 0.15
       WIDTH 1.50 PARALLEL 1.5 WITHIN 0.50 LONGJOGSPACING 0.30 ; " ;

    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 ;
        SPACING 0.080 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ;
        SPACING 0.100 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ENCLOSECUT BELOW 0.050 CUTSPACING 0.145 ALLCUTS ;" ;

    #MxLPC: Cap Rule 
    PROPERTY LEF58_SPACING "
	SPACING 0.115 ENDOFLINE 0.055 WITHIN 0.000 PARALLELEDGE 0.060 WITHIN 0.120 MINLENGTH 0.150 TWOEDGES SAMEMETAL ; " ;

#    #  BR.S1 BR.S2 BR.S3  #
#    PROPERTY LEF58_SPACING "
#      SPACING 0.236 CONVEXCORNERS EXTENSION 0.16 0.23 ;
#      SPACING 0.080 CONVEXCORNERS EXTENSION 0.23 0.075 SINGLE 0.3 0.08 0.12 SPANLENGTH 0.3 OPPOSITEWIDTH 0.055 OPPOSITEEXTENSION 0.055 0.025 0.1 ;
#      SPACING 0.051 CONVEXCORNERS EXTENSION 0.160 0.115 SAMESIDE 0.09 ; " ;

    

    PROPERTY LEF58_MINIMUMCUT "    
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 WITHIN 0.100000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 4 CUTCLASS VDOUBLECUT 2 WIDTH 0.440000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000  LENGTH 0.180000 WITHIN 1.651000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.000000  LENGTH 1.000000 WITHIN 4.001000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.500000  LENGTH 5.000000 WITHIN 10.001000 ; " ; 

    HEIGHT 0.465 ;
    THICKNESS 0.090000 ;
    FILLACTIVESPACING 0.2 ;
    RESISTANCE RPERSQ 0.428 ;
    CAPACITANCE CPERSQDIST 0.000312857 ;
    EDGECAPACITANCE 7.44E-05 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 9.123323 8.283339 7.737038 7.736060 6.463440 6.055773 5.823409 5.684512 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 32.681533 33.848730 34.237219 17.118898 17.391244 17.449604 17.478784 17.494995 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

END M2

LAYER VIA2
    TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
        CUTCLASS VSINGLECUT WIDTH 0.05 LENGTH 0.05 CUTS 1 ;
        CUTCLASS VDOUBLECUT WIDTH 0.05 LENGTH 0.13 CUTS 2 ;" ;

    #EFP.VIAx.S.1~6
    PROPERTY LEF58_EOLSPACING "
        EOLSPACING 0.08 0.09 CUTCLASS VSINGLECUT TO VDOUBLECUT 0.085 0.09 ENDWIDTH 0.07 PRL -0.04
        ENCLOSURE 0.04 0.00 EXTENSION 0.065 0.12 SPANLENGTH 0.055 ; " ;

    PROPERTY LEF58_SPACINGTABLE "
    	SPACINGTABLE PRL -0.04 MAXXY 
    	CUTCLASS	VSINGLECUT	VDOUBLECUT
    	VSINGLECUT	0.070 0.080	0.075 0.080
    	VDOUBLECUT	0.075 0.080	0.080 0.080 ;" ;

    #Enhanced Mx.S.8
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VSINGLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VDOUBLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;

    #VIAx.R.10R
    PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE LAYER VIA1 PRL 0.02
      CUTCLASS    VSINGLECUT  VDOUBLECUT
      VSINGLECUT  0.000 0.060 0.000 0.060
      VDOUBLECUT  0.000 0.060 0.000 0.060 ;" ;

    
    PROPERTY LEF58_ENCLOSUREEDGE "
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ; 
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1  ;
        ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1 ; " ;
        
 
    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS VSINGLECUT 0 0.03 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.02 0.02 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.01 0.025 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.02 SIDE 0.02 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.03 SIDE 0.01 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.01 SIDE 0.03 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.04 SIDE 0 ;
        " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ;
    DCCURRENTDENSITY	AVERAGE
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ; 

END VIA2

LAYER M3
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.100 0.100 ;
    OFFSET 0.000 0.000 ;
    MINWIDTH 0.050000 ;
    MAXWIDTH 4.500000 ;
    WIDTH 0.050000 ;

    AREA 0.017 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.050000 MAXEDGES 1 ;
    PROPERTY LEF58_MINSTEP "MINSTEP 0.05 MAXEDGES 1 MINADJACENTLENGTH 0.065 CONVEXCORNER ;" ;
    PROPERTY LEF58_AREA "AREA 0.044000 EXCEPTEDGELENGTH 0.130000 EXCEPTMINSIZE 0.050000 0.130000 ;" ;

    #---RR:RE:EFP.Mx.S.3 hook v01---#
    SPACING 0.07 NOTCHLENGTH 0.155 ;


    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.220000  0.470000  0.630000  1.500000
      WIDTH  0.000000  0.050000  0.050000  0.050000  0.050000  0.050000
      WIDTH  0.090000  0.050000  0.060000  0.060000  0.060000  0.060000
      WIDTH  0.130000  0.050000  0.080000  0.080000  0.080000  0.080000
      WIDTH  0.160000  0.050000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.470000  0.050000  0.100000  0.130000  0.130000  0.130000
      WIDTH  0.630000  0.050000  0.100000  0.130000  0.150000  0.150000
      WIDTH  1.500000  0.050000  0.100000  0.130000  0.150000  0.500000 ;
    
    PROPERTY LEF58_SPACINGTABLE "
       SPACINGTABLE JOGTOJOGSPACING 0.3 JOGWIDTH 0.22
       SHORTJOGSPACING 0.06
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.29 LONGJOGSPACING 0.08
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.19 LONGJOGSPACING 0.10
       WIDTH 0.47 PARALLEL 0.5 WITHIN 0.32 LONGJOGSPACING 0.13
       WIDTH 0.63 PARALLEL 0.7 WITHIN 0.34 LONGJOGSPACING 0.15
       WIDTH 1.50 PARALLEL 1.5 WITHIN 0.50 LONGJOGSPACING 0.30 ; " ;

    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 ;
        SPACING 0.080 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ;
        SPACING 0.100 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ENCLOSECUT BELOW 0.050 CUTSPACING 0.145 ALLCUTS ;" ;

    #MxLPC: Cap Rule 
    PROPERTY LEF58_SPACING "
	SPACING 0.115 ENDOFLINE 0.055 WITHIN 0.000 PARALLELEDGE 0.060 WITHIN 0.120 MINLENGTH 0.150 TWOEDGES SAMEMETAL ; " ;

#    #  BR.S1 BR.S2 BR.S3  #
#    PROPERTY LEF58_SPACING "
#      SPACING 0.236 CONVEXCORNERS EXTENSION 0.16 0.23 ;
#      SPACING 0.080 CONVEXCORNERS EXTENSION 0.23 0.075 SINGLE 0.3 0.08 0.12 SPANLENGTH 0.3 OPPOSITEWIDTH 0.055 OPPOSITEEXTENSION 0.055 0.025 0.1 ;
#      SPACING 0.051 CONVEXCORNERS EXTENSION 0.160 0.115 SAMESIDE 0.09 ; " ;

    #Mx_S_37R
    PROPERTY LEF58_CORNERFILLSPACING "CORNERFILLSPACING 0.05 EDGELENGTH 0.05 0.12  ADJACENTEOL 0.06 ;" ;


    PROPERTY LEF58_MINIMUMCUT "    
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 WITHIN 0.100000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 4 CUTCLASS VDOUBLECUT 2 WIDTH 0.440000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000  LENGTH 0.180000 WITHIN 1.651000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.000000  LENGTH 1.000000 WITHIN 4.001000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.500000  LENGTH 5.000000 WITHIN 10.001000 ; " ; 

    HEIGHT 0.565 ;
    THICKNESS 0.090000 ;
    FILLACTIVESPACING 0.2 ;
    RESISTANCE RPERSQ 0.428 ;
    CAPACITANCE CPERSQDIST 0.000312857 ;
    EDGECAPACITANCE 7.44E-05 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 8.832119 7.803326 7.134792 7.133588 5.521506 4.975651 4.654273 4.457723 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 32.681533 33.848730 34.237219 17.118898 17.391244 17.449604 17.478784 17.494995 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

END M3

LAYER VIA3
    TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
        CUTCLASS VSINGLECUT WIDTH 0.05 LENGTH 0.05 CUTS 1 ;
        CUTCLASS VDOUBLECUT WIDTH 0.05 LENGTH 0.13 CUTS 2 ;" ;

    #EFP.VIAx.S.1~6
    PROPERTY LEF58_EOLSPACING "
        EOLSPACING 0.08 0.09 CUTCLASS VSINGLECUT TO VDOUBLECUT 0.085 0.09 ENDWIDTH 0.07 PRL -0.04
        ENCLOSURE 0.04 0.00 EXTENSION 0.065 0.12 SPANLENGTH 0.055 ; " ;

    PROPERTY LEF58_SPACINGTABLE "
    	SPACINGTABLE PRL -0.04 MAXXY 
    	CUTCLASS	VSINGLECUT	VDOUBLECUT
    	VSINGLECUT	0.070 0.080	0.075 0.080
    	VDOUBLECUT	0.075 0.080	0.080 0.080 ;" ;

    #Enhanced Mx.S.8
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VSINGLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VDOUBLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;

    #VIAx.R.10R
    PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE LAYER VIA2 PRL 0.02
      CUTCLASS    VSINGLECUT  VDOUBLECUT
      VSINGLECUT  0.000 0.060 0.000 0.060
      VDOUBLECUT  0.000 0.060 0.000 0.060 ;" ;

    
    PROPERTY LEF58_ENCLOSUREEDGE "
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ; 
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1  ;
        ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1 ; " ;
        
 
    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS VSINGLECUT 0 0.03 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.02 0.02 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.01 0.025 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.02 SIDE 0.02 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.03 SIDE 0.01 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.01 SIDE 0.03 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.04 SIDE 0 ;
        " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ;
    DCCURRENTDENSITY	AVERAGE
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ; 

END VIA3

LAYER M4
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.100 0.100 ;
    OFFSET 0.000 0.000 ;
    MINWIDTH 0.050000 ;
    MAXWIDTH 4.500000 ;
    WIDTH 0.050000 ;

    AREA 0.017 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.050000 MAXEDGES 1 ;
    PROPERTY LEF58_MINSTEP "MINSTEP 0.05 MAXEDGES 1 MINADJACENTLENGTH 0.065 CONVEXCORNER ;" ;
    PROPERTY LEF58_AREA "AREA 0.044000 EXCEPTEDGELENGTH 0.130000 EXCEPTMINSIZE 0.050000 0.130000 ;" ;

    #---RR:RE:EFP.Mx.S.3 hook v01---#
    SPACING 0.07 NOTCHLENGTH 0.155 ;


    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.220000  0.470000  0.630000  1.500000
      WIDTH  0.000000  0.050000  0.050000  0.050000  0.050000  0.050000
      WIDTH  0.090000  0.050000  0.060000  0.060000  0.060000  0.060000
      WIDTH  0.130000  0.050000  0.080000  0.080000  0.080000  0.080000
      WIDTH  0.160000  0.050000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.470000  0.050000  0.100000  0.130000  0.130000  0.130000
      WIDTH  0.630000  0.050000  0.100000  0.130000  0.150000  0.150000
      WIDTH  1.500000  0.050000  0.100000  0.130000  0.150000  0.500000 ;
    
    PROPERTY LEF58_SPACINGTABLE "
       SPACINGTABLE JOGTOJOGSPACING 0.3 JOGWIDTH 0.22
       SHORTJOGSPACING 0.06
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.29 LONGJOGSPACING 0.08
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.19 LONGJOGSPACING 0.10
       WIDTH 0.47 PARALLEL 0.5 WITHIN 0.32 LONGJOGSPACING 0.13
       WIDTH 0.63 PARALLEL 0.7 WITHIN 0.34 LONGJOGSPACING 0.15
       WIDTH 1.50 PARALLEL 1.5 WITHIN 0.50 LONGJOGSPACING 0.30 ; " ;

    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 ;
        SPACING 0.080 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ;
        SPACING 0.100 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ENCLOSECUT BELOW 0.050 CUTSPACING 0.145 ALLCUTS ;" ;

    #MxLPC: Cap Rule 
    PROPERTY LEF58_SPACING "
	SPACING 0.115 ENDOFLINE 0.055 WITHIN 0.000 PARALLELEDGE 0.060 WITHIN 0.120 MINLENGTH 0.150 TWOEDGES SAMEMETAL ; " ;

#    #  BR.S1 BR.S2 BR.S3  #
#    PROPERTY LEF58_SPACING "
#      SPACING 0.236 CONVEXCORNERS EXTENSION 0.16 0.23 ;
#      SPACING 0.080 CONVEXCORNERS EXTENSION 0.23 0.075 SINGLE 0.3 0.08 0.12 SPANLENGTH 0.3 OPPOSITEWIDTH 0.055 OPPOSITEEXTENSION 0.055 0.025 0.1 ;
#      SPACING 0.051 CONVEXCORNERS EXTENSION 0.160 0.115 SAMESIDE 0.09 ; " ;

    #Mx_S_37R
    PROPERTY LEF58_CORNERFILLSPACING "CORNERFILLSPACING 0.05 EDGELENGTH 0.05 0.12  ADJACENTEOL 0.06 ;" ;


    PROPERTY LEF58_MINIMUMCUT "    
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 WITHIN 0.100000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 4 CUTCLASS VDOUBLECUT 2 WIDTH 0.440000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000  LENGTH 0.180000 WITHIN 1.651000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.000000  LENGTH 1.000000 WITHIN 4.001000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.500000  LENGTH 5.000000 WITHIN 10.001000 ; " ; 

    HEIGHT 0.665 ;
    THICKNESS 0.090000 ;
    FILLACTIVESPACING 0.2 ;
    RESISTANCE RPERSQ 0.428 ;
    CAPACITANCE CPERSQDIST 0.000312857 ;
    EDGECAPACITANCE 7.44E-05 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 8.695460 7.582195 6.856247 6.854934 5.065452 4.436161 4.056050 3.818898 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 32.681533 33.848730 34.237219 17.118898 17.391244 17.449604 17.478784 17.494995 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

END M4

LAYER VIA4
    TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
        CUTCLASS VSINGLECUT WIDTH 0.05 LENGTH 0.05 CUTS 1 ;
        CUTCLASS VDOUBLECUT WIDTH 0.05 LENGTH 0.13 CUTS 2 ;" ;

    #EFP.VIAx.S.1~6
    PROPERTY LEF58_EOLSPACING "
        EOLSPACING 0.08 0.09 CUTCLASS VSINGLECUT TO VDOUBLECUT 0.085 0.09 ENDWIDTH 0.07 PRL -0.04
        ENCLOSURE 0.04 0.00 EXTENSION 0.065 0.12 SPANLENGTH 0.055 ; " ;

    PROPERTY LEF58_SPACINGTABLE "
    	SPACINGTABLE PRL -0.04 MAXXY 
    	CUTCLASS	VSINGLECUT	VDOUBLECUT
    	VSINGLECUT	0.070 0.080	0.075 0.080
    	VDOUBLECUT	0.075 0.080	0.080 0.080 ;" ;

    #Enhanced Mx.S.8
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VSINGLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VDOUBLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;

    #VIAx.R.10R
    PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE LAYER VIA3 PRL 0.02
      CUTCLASS    VSINGLECUT  VDOUBLECUT
      VSINGLECUT  0.000 0.060 0.000 0.060
      VDOUBLECUT  0.000 0.060 0.000 0.060 ;" ;

    
    PROPERTY LEF58_ENCLOSUREEDGE "
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ; 
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1  ;
        ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1 ; " ;
        
 
    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS VSINGLECUT 0 0.03 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.02 0.02 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.01 0.025 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.02 SIDE 0.02 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.03 SIDE 0.01 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.01 SIDE 0.03 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.04 SIDE 0 ;
        " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ;
    DCCURRENTDENSITY	AVERAGE
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ; 

END VIA4

LAYER M5
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.100 0.100 ;
    OFFSET 0.000 0.000 ;
    MINWIDTH 0.050000 ;
    MAXWIDTH 4.500000 ;
    WIDTH 0.050000 ;

    AREA 0.017 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.050000 MAXEDGES 1 ;
    PROPERTY LEF58_MINSTEP "MINSTEP 0.05 MAXEDGES 1 MINADJACENTLENGTH 0.065 CONVEXCORNER ;" ;
    PROPERTY LEF58_AREA "AREA 0.044000 EXCEPTEDGELENGTH 0.130000 EXCEPTMINSIZE 0.050000 0.130000 ;" ;

    #---RR:RE:EFP.Mx.S.3 hook v01---#
    SPACING 0.07 NOTCHLENGTH 0.155 ;


    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.220000  0.470000  0.630000  1.500000
      WIDTH  0.000000  0.050000  0.050000  0.050000  0.050000  0.050000
      WIDTH  0.090000  0.050000  0.060000  0.060000  0.060000  0.060000
      WIDTH  0.130000  0.050000  0.080000  0.080000  0.080000  0.080000
      WIDTH  0.160000  0.050000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.470000  0.050000  0.100000  0.130000  0.130000  0.130000
      WIDTH  0.630000  0.050000  0.100000  0.130000  0.150000  0.150000
      WIDTH  1.500000  0.050000  0.100000  0.130000  0.150000  0.500000 ;
    
    PROPERTY LEF58_SPACINGTABLE "
       SPACINGTABLE JOGTOJOGSPACING 0.3 JOGWIDTH 0.22
       SHORTJOGSPACING 0.06
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.29 LONGJOGSPACING 0.08
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.19 LONGJOGSPACING 0.10
       WIDTH 0.47 PARALLEL 0.5 WITHIN 0.32 LONGJOGSPACING 0.13
       WIDTH 0.63 PARALLEL 0.7 WITHIN 0.34 LONGJOGSPACING 0.15
       WIDTH 1.50 PARALLEL 1.5 WITHIN 0.50 LONGJOGSPACING 0.30 ; " ;

    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 ;
        SPACING 0.080 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ;
        SPACING 0.100 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ENCLOSECUT BELOW 0.050 CUTSPACING 0.145 ALLCUTS ;" ;

    #MxLPC: Cap Rule 
    PROPERTY LEF58_SPACING "
	SPACING 0.115 ENDOFLINE 0.055 WITHIN 0.000 PARALLELEDGE 0.060 WITHIN 0.120 MINLENGTH 0.150 TWOEDGES SAMEMETAL ; " ;

#    #  BR.S1 BR.S2 BR.S3  #
#    PROPERTY LEF58_SPACING "
#      SPACING 0.236 CONVEXCORNERS EXTENSION 0.16 0.23 ;
#      SPACING 0.080 CONVEXCORNERS EXTENSION 0.23 0.075 SINGLE 0.3 0.08 0.12 SPANLENGTH 0.3 OPPOSITEWIDTH 0.055 OPPOSITEEXTENSION 0.055 0.025 0.1 ;
#      SPACING 0.051 CONVEXCORNERS EXTENSION 0.160 0.115 SAMESIDE 0.09 ; " ;

    #Mx_S_37R
    PROPERTY LEF58_CORNERFILLSPACING "CORNERFILLSPACING 0.05 EDGELENGTH 0.05 0.12  ADJACENTEOL 0.06 ;" ;


    PROPERTY LEF58_MINIMUMCUT "    
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 WITHIN 0.100000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 4 CUTCLASS VDOUBLECUT 2 WIDTH 0.440000  ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000  LENGTH 0.180000 WITHIN 1.651000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.000000  LENGTH 1.000000 WITHIN 4.001000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.500000  LENGTH 5.000000 WITHIN 10.001000 ; " ; 

    HEIGHT 0.765 ;
    THICKNESS 0.090000 ;
    FILLACTIVESPACING 0.2 ;
    RESISTANCE RPERSQ 0.428 ;
    CAPACITANCE CPERSQDIST 0.000312857 ;
    EDGECAPACITANCE 7.44E-05 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 8.636347 7.472521 6.711398 6.710018 4.805843 4.117744 3.693471 3.424119 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 32.681533 33.848730 34.237219 17.118898 17.391244 17.449604 17.478784 17.494995 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

END M5

LAYER VIA5
    TYPE CUT ;

    PROPERTY LEF58_CUTCLASS "
        CUTCLASS VSINGLECUT WIDTH 0.05 LENGTH 0.05 CUTS 1 ;
        CUTCLASS VDOUBLECUT WIDTH 0.05 LENGTH 0.13 CUTS 2 ;" ;

    #EFP.VIAx.S.1~6
    PROPERTY LEF58_EOLSPACING "
        EOLSPACING 0.08 0.09 CUTCLASS VSINGLECUT TO VDOUBLECUT 0.085 0.09 ENDWIDTH 0.07 PRL -0.04
        ENCLOSURE 0.04 0.00 EXTENSION 0.065 0.12 SPANLENGTH 0.055 ; " ;

    PROPERTY LEF58_SPACINGTABLE "
    	SPACINGTABLE PRL -0.04 MAXXY 
    	CUTCLASS	VSINGLECUT	VDOUBLECUT
    	VSINGLECUT	0.070 0.080	0.075 0.080
    	VDOUBLECUT	0.075 0.080	0.080 0.080 ;" ;

    #Enhanced Mx.S.8
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VSINGLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;
    PROPERTY LEF58_EOLENCLOSURE "
        EOLENCLOSURE 0.070 CUTCLASS VDOUBLECUT ABOVE 0.030 PARALLELEDGE 0.115 EXTENSION 0.070 0.025 MINLENGTH 0.050 ; " ;

    #VIAx.R.10R
    PROPERTY LEF58_SPACINGTABLE "
      SPACINGTABLE LAYER VIA4 PRL 0.02
      CUTCLASS    VSINGLECUT  VDOUBLECUT
      VSINGLECUT  0.000 0.060 0.000 0.060
      VDOUBLECUT  0.000 0.060 0.000 0.060 ;" ;

    
    PROPERTY LEF58_ENCLOSUREEDGE "
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ; 
    	ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT 0.015000 WIDTH 0.160500 PARALLEL 0.100000 WITHIN 0.130000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.010000 WIDTH 0.070500 PARALLEL 0.100000 WITHIN 0.100000 ;
    	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.055500 PARALLEL 0.100000 WITHIN 0.065000 ;
	ENCLOSUREEDGE CUTCLASS VDOUBLECUT  0.005000 WIDTH 0.050500 PARALLEL 0.100000 WITHIN 0.060000 EXCEPTTWOEDGES ;
        ENCLOSUREEDGE CUTCLASS VSINGLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1  ;
        ENCLOSUREEDGE CUTCLASS VDOUBLECUT ABOVE 0.01 CONVEXCORNERS 0.120 0.060 PARALLEL 0.051 LENGTH 0.1 ; " ;
        
 
    PROPERTY LEF58_ENCLOSURE "
        ENCLOSURE CUTCLASS VSINGLECUT 0 0.03 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.02 0.02 ;
        ENCLOSURE CUTCLASS VSINGLECUT 0.01 0.025 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.02 SIDE 0.02 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.03 SIDE 0.01 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.01 SIDE 0.03 ;
        ENCLOSURE CUTCLASS VDOUBLECUT END 0.04 SIDE 0 ;
        " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ;
    DCCURRENTDENSITY	AVERAGE
        CUTAREA         0.0025 0.0065 ;
        TABLEENTRIES	20.641975 15.878443 ; 

END VIA5

LAYER M6
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.100 0.100 ;
    OFFSET 0.000 0.000 ;
    MINWIDTH 0.050000 ;
    MAXWIDTH 4.500000 ;
    WIDTH 0.050000 ;

    AREA 0.017 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.050000 MAXEDGES 1 ;
    PROPERTY LEF58_MINSTEP "MINSTEP 0.05 MAXEDGES 1 MINADJACENTLENGTH 0.065 CONVEXCORNER ;" ;
    PROPERTY LEF58_AREA "AREA 0.044000 EXCEPTEDGELENGTH 0.130000 EXCEPTMINSIZE 0.050000 0.130000 ;" ;

    #---RR:RE:EFP.Mx.S.3 hook v01---#
    SPACING 0.07 NOTCHLENGTH 0.155 ;


    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.220000  0.470000  0.630000  1.500000
      WIDTH  0.000000  0.050000  0.050000  0.050000  0.050000  0.050000
      WIDTH  0.090000  0.050000  0.060000  0.060000  0.060000  0.060000
      WIDTH  0.130000  0.050000  0.080000  0.080000  0.080000  0.080000
      WIDTH  0.160000  0.050000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.470000  0.050000  0.100000  0.130000  0.130000  0.130000
      WIDTH  0.630000  0.050000  0.100000  0.130000  0.150000  0.150000
      WIDTH  1.500000  0.050000  0.100000  0.130000  0.150000  0.500000 ;
    
    PROPERTY LEF58_SPACINGTABLE "
       SPACINGTABLE JOGTOJOGSPACING 0.3 JOGWIDTH 0.22
       SHORTJOGSPACING 0.06
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.29 LONGJOGSPACING 0.08
       WIDTH 0.25 PARALLEL 0.3 WITHIN 0.19 LONGJOGSPACING 0.10
       WIDTH 0.47 PARALLEL 0.5 WITHIN 0.32 LONGJOGSPACING 0.13
       WIDTH 0.63 PARALLEL 0.7 WITHIN 0.34 LONGJOGSPACING 0.15
       WIDTH 1.50 PARALLEL 1.5 WITHIN 0.50 LONGJOGSPACING 0.30 ; " ;

    PROPERTY LEF58_SPACING "
        SPACING 0.070 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 ;
        SPACING 0.080 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ;
        SPACING 0.100 ENDOFLINE 0.070 WITHIN 0.025 ENDTOEND 0.080 PARALLELEDGE SUBTRACTEOLWIDTH 0.115 WITHIN 0.070 MINLENGTH 0.050 ENCLOSECUT BELOW 0.050 CUTSPACING 0.145 ALLCUTS ;" ;

    #MxLPC: Cap Rule 
    PROPERTY LEF58_SPACING "
	SPACING 0.115 ENDOFLINE 0.055 WITHIN 0.000 PARALLELEDGE 0.060 WITHIN 0.120 MINLENGTH 0.150 TWOEDGES SAMEMETAL ; " ;

#    #  BR.S1 BR.S2 BR.S3  #
#    PROPERTY LEF58_SPACING "
#      SPACING 0.236 CONVEXCORNERS EXTENSION 0.16 0.23 ;
#      SPACING 0.080 CONVEXCORNERS EXTENSION 0.23 0.075 SINGLE 0.3 0.08 0.12 SPANLENGTH 0.3 OPPOSITEWIDTH 0.055 OPPOSITEEXTENSION 0.055 0.025 0.1 ;
#      SPACING 0.051 CONVEXCORNERS EXTENSION 0.160 0.115 SAMESIDE 0.09 ; " ;

    #Mx_S_37R
    PROPERTY LEF58_CORNERFILLSPACING "CORNERFILLSPACING 0.05 EDGELENGTH 0.05 0.12  ADJACENTEOL 0.06 ;" ;


    PROPERTY LEF58_MINIMUMCUT "    
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 WITHIN 0.100000 FROMBELOW ;
    MINIMUMCUT CUTCLASS VSINGLECUT 4 CUTCLASS VDOUBLECUT 2 WIDTH 0.440000 FROMBELOW ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 0.180000 FROMBELOW LENGTH 0.180000 WITHIN 1.651000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.000000 FROMBELOW LENGTH 1.000000 WITHIN 4.001000 ;
    MINIMUMCUT CUTCLASS VSINGLECUT 2 CUTCLASS VDOUBLECUT 1 WIDTH 1.500000 FROMBELOW LENGTH 5.000000 WITHIN 10.001000 ;
    MINIMUMCUT 2 WIDTH 0.300000 FROMABOVE ;
    MINIMUMCUT 4 WIDTH 0.700000 FROMABOVE ;
    MINIMUMCUT 2 WIDTH 0.300000 FROMABOVE LENGTH 0.300000 WITHIN 0.801000 ;
    MINIMUMCUT 2 WIDTH 2.000000 FROMABOVE LENGTH 2.000000 WITHIN 2.001000 ;
    MINIMUMCUT 2 WIDTH 3.000000 FROMABOVE LENGTH 10.000000 WITHIN 5.001000 ; " ; 

    HEIGHT 0.865 ;
    THICKNESS 0.090000 ;
    FILLACTIVESPACING 0.2 ;
    RESISTANCE RPERSQ 0.428 ;
    CAPACITANCE CPERSQDIST 0.000312857 ;
    EDGECAPACITANCE 7.44E-05 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 8.596164 7.399856 6.615760 6.614335 4.631802 3.900541 3.441973 3.146355 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 32.681533 33.848730 34.237219 17.118898 17.391244 17.449604 17.478784 17.494995 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.045000 0.090000 0.134900 0.135000 0.450000 0.900000 1.800000 4.050000 ;
        TABLEENTRIES	 0.929600 0.962800 0.973850 0.973867 0.989360 0.992680 0.994340 0.995262 ;

END M6

LAYER VIA6
    TYPE CUT ;
    SPACING 0.100000 ;
    SPACING 0.130000 ADJACENTCUTS 3 WITHIN 0.140000 ;

    PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ; " ;

    ENCLOSURE BELOW 0.015 0.04 ;
    ENCLOSURE ABOVE 0 0.04 ;
    ENCLOSURE ABOVE 0.03 0.03 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	20.172840 ;
    DCCURRENTDENSITY	AVERAGE 20.172840 ; 

END VIA6

LAYER M7
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.200000 0.200000 ;
    OFFSET 0.000000 0.000000 ;
    MINWIDTH 0.100000 ;
    MAXWIDTH 12.000000 ;
    WIDTH 0.100000 ;

    AREA 0.052000 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.100000 MAXEDGES 1 ;

    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.380000  0.400000  1.500000  4.500000
      WIDTH  0.000000  0.100000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.200000  0.100000  0.120000  0.120000  0.120000  0.120000
      WIDTH  0.400000  0.100000  0.120000  0.160000  0.160000  0.160000
      WIDTH  1.500000  0.100000  0.120000  0.160000  0.500000  0.500000
      WIDTH  4.500000  0.100000  0.120000  0.160000  0.500000  1.500000 ;

    
    MINIMUMCUT 2 WIDTH 0.300000  ;
    MINIMUMCUT 4 WIDTH 0.700000  ;
    MINIMUMCUT 2 WIDTH 0.300000  LENGTH 0.300000 WITHIN 0.801000 ;
    MINIMUMCUT 2 WIDTH 2.000000  LENGTH 2.000000 WITHIN 2.001000 ;
    MINIMUMCUT 2 WIDTH 3.000000  LENGTH 10.000000 WITHIN 5.001000 ;

    HEIGHT 0.965 ;
    THICKNESS 0.190000 ;
    FILLACTIVESPACING 0.3 ;

    PROPERTY LEF58_SPACING "SPACING 0.120 ENDOFLINE 0.120 WITHIN 0.035 PARALLELEDGE 0.120 WITHIN 0.120 MINLENGTH 0.100 ; " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 1.815467 1.946117 1.946311 2.129493 2.168747 2.189406 2.201458 2.204729 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 9.451966 8.777560 8.776081 6.246066 5.157677 4.395805 3.850152 3.683622 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 30.814142 33.031689 16.517491 18.072078 18.405204 18.580533 18.682809 18.710569 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 1.815467 1.946117 1.946311 2.129493 2.168747 2.189406 2.201458 2.204729 ;

    RESISTANCE RPERSQ	0.4280000000 ;
    CAPACITANCE CPERSQDIST	0.0004911111 ;
    EDGECAPACITANCE	0.0000674000 ;
END M7

LAYER VIA7
    TYPE CUT ;
    SPACING 0.100000 ;
    SPACING 0.130000 ADJACENTCUTS 3 WITHIN 0.140000 ;

    PROPERTY LEF58_SPACING "SPACING 0.13 PARALLELOVERLAP EXCEPTSAMENET ; " ;

    ENCLOSURE BELOW 0 0.04 ;
    ENCLOSURE ABOVE 0 0.04 ;
    ENCLOSURE  0.03 0.03 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	20.172840 ;
    DCCURRENTDENSITY	AVERAGE 20.172840 ; 

END VIA7

LAYER M8
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.200000 0.200000 ;
    OFFSET 0.000000 0.000000 ;
    MINWIDTH 0.100000 ;
    MAXWIDTH 12.000000 ;
    WIDTH 0.100000 ;

    AREA 0.052000 ;
    MINENCLOSEDAREA 0.200000 ;
    MINSTEP 0.100000 MAXEDGES 1 ;

    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  0.380000  0.400000  1.500000  4.500000
      WIDTH  0.000000  0.100000  0.100000  0.100000  0.100000  0.100000
      WIDTH  0.200000  0.100000  0.120000  0.120000  0.120000  0.120000
      WIDTH  0.400000  0.100000  0.120000  0.160000  0.160000  0.160000
      WIDTH  1.500000  0.100000  0.120000  0.160000  0.500000  0.500000
      WIDTH  4.500000  0.100000  0.120000  0.160000  0.500000  1.500000 ;

    
    MINIMUMCUT 2 WIDTH 0.300000 FROMBELOW ;
    MINIMUMCUT 4 WIDTH 0.700000 FROMBELOW ;
    MINIMUMCUT 2 WIDTH 0.300000 FROMBELOW LENGTH 0.300000 WITHIN 0.801000 ;
    MINIMUMCUT 2 WIDTH 2.000000 FROMBELOW LENGTH 2.000000 WITHIN 2.001000 ;
    MINIMUMCUT 2 WIDTH 3.000000 FROMBELOW LENGTH 10.000000 WITHIN 5.001000 ;
    MINIMUMCUT 2 WIDTH 1.800000 FROMABOVE ;
    MINIMUMCUT 2 WIDTH 3.000000 FROMABOVE LENGTH 10.000000 WITHIN 5.001000 ; 

    HEIGHT 1.175 ;
    THICKNESS 0.190000 ;
    FILLACTIVESPACING 0.3 ;

    PROPERTY LEF58_SPACING "SPACING 0.120 ENDOFLINE 0.120 WITHIN 0.035 PARALLELEDGE 0.120 WITHIN 0.120 MINLENGTH 0.100 ; " ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 1.815467 1.946117 1.946311 2.129493 2.168747 2.189406 2.201458 2.204729 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 9.391159 8.696031 8.694511 6.089599 4.953915 4.146139 3.556351 3.373587 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 30.814142 33.031689 16.517491 18.072078 18.405204 18.580533 18.682809 18.710569 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.090000 0.134900 0.135000 0.450000 0.900000 1.900000 5.400000 10.800000 ;
        TABLEENTRIES	 1.815467 1.946117 1.946311 2.129493 2.168747 2.189406 2.201458 2.204729 ;

    RESISTANCE RPERSQ	0.4280000000 ;
    CAPACITANCE CPERSQDIST	0.0004911111 ;
    EDGECAPACITANCE	0.0000674000 ;
END M8

LAYER VIA8
    TYPE CUT ;
    SPACING 0.340000 ;
    SPACING 0.540000 ADJACENTCUTS 3 WITHIN 0.560000 ;

    ENCLOSURE 0.02 0.08 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	20.486587 ;
    DCCURRENTDENSITY	AVERAGE 20.486587 ; 

END VIA8

LAYER M9
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH 0.800000 0.800000 ;
    OFFSET 0.000000 0.000000 ;
    MINWIDTH 0.400000 ;
    MAXWIDTH 12.000000 ;
    WIDTH 0.400000 ;

    AREA 0.565000 ;
    MINENCLOSEDAREA 0.565000 ;

    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  1.500000  4.500000
      WIDTH  0.000000  0.400000  0.400000  0.400000
      WIDTH  1.500000  0.400000  0.500000  0.500000
      WIDTH  4.500000  0.400000  0.500000  1.500000 ;

    
    MINIMUMCUT 2 WIDTH 1.800000  ;
    MINIMUMCUT 2 WIDTH 3.000000  LENGTH 10.000000 WITHIN 5.001000 ; 

    HEIGHT 1.385 ;
    THICKNESS 0.850000 ;
    FILLACTIVESPACING 0.6 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 43000.011 ) ( 0.2 43091.2 ) ( 0.5 43228.0 ) ( 1 43456 ) ( 1.5 43684.0 ) ) ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 8.545333 8.846933 8.947467 8.997733 9.022867 9.031244 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 13.511040 10.129349 8.457550 7.422844 6.830258 6.618339 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 77.601041 80.339901 81.252855 81.709331 81.937570 82.013649 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 8.545333 8.846933 8.947467 8.997733 9.022867 9.031244 ;

    RESISTANCE RPERSQ 0.022 ;
    CAPACITANCE CPERSQDIST 6.025E-05 ;
    EDGECAPACITANCE 9.3E-05 ;
END M9

LAYER VIA9
    TYPE CUT ;
    SPACING 0.340000 ;
    SPACING 0.540000 ADJACENTCUTS 3 WITHIN 0.560000 ;

    ENCLOSURE 0.02 0.08 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 900 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 99999 ) ( 0.2 99999 ) ( 0.5 99999 ) ) ;
    ANTENNACUMDIFFAREARATIO PWL ( ( 0 50 ) ( 0.000025 900.00525 ) ( 0.2 942.0 ) ( 0.5 1005.0 ) ( 1 1110 ) ( 1.5 1215.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	29.311462 ;
    DCCURRENTDENSITY	AVERAGE 29.311462 ; 

END VIA9

LAYER M10
    TYPE ROUTING ;
    DIRECTION HORIZONTAL ;
    PITCH 0.800000 0.800000 ;
    OFFSET 0.000000 0.000000 ;
    MINWIDTH 0.400000 ;
    MAXWIDTH 12.000000 ;
    WIDTH 0.400000 ;

    AREA 0.565000 ;
    MINENCLOSEDAREA 0.565000 ;

    SPACINGTABLE
    PARALLELRUNLENGTH  0.000000  1.500000  4.500000
      WIDTH  0.000000  0.400000  0.400000  0.400000
      WIDTH  1.500000  0.400000  0.500000  0.500000
      WIDTH  4.500000  0.400000  0.500000  1.500000 ;

    
    MINIMUMCUT 2 WIDTH 1.800000 FROMBELOW ;
    MINIMUMCUT 2 WIDTH 3.000000 FROMBELOW LENGTH 10.000000 WITHIN 5.001000 ; 

    HEIGHT 2.245 ;
    THICKNESS 0.850000 ;
    FILLACTIVESPACING 0.6 ;

    
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 5000 ) ( 0.000025 50000.2 ) ( 0.2 51600.0 ) ( 0.5 54000.0 ) ( 1 58000 ) ( 1.5 62000.0 ) ) ;
    ANTENNACUMAREARATIO 5000 ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 1000 ) ( 0.000025 50000.2 ) ( 0.2 51600.0 ) ( 0.5 54000.0 ) ( 1 58000 ) ( 1.5 62000.0 ) ) ;
    ANTENNACUMAREARATIO 1000 ;

    MINIMUMDENSITY      10 ;
    MAXIMUMDENSITY      85 ;
    DENSITYCHECKWINDOW 125 125 ;
    DENSITYCHECKSTEP    62.5 ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 8.545333 8.846933 8.947467 8.997733 9.022867 9.031244 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 13.326086 9.843819 8.096877 6.999265 6.361867 6.131865 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 77.601041 80.339901 81.252855 81.709331 81.937570 82.013649 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 0.360000 0.900000 1.800000 3.600000 7.200000 10.800000 ;
        TABLEENTRIES	 8.545333 8.846933 8.947467 8.997733 9.022867 9.031244 ;

    RESISTANCE RPERSQ 0.022 ;
    CAPACITANCE CPERSQDIST 6.025E-05 ;
    EDGECAPACITANCE 9.3E-05 ;
END M10

LAYER RV
    TYPE CUT ;
    SPACING 2.00 ;

    ENCLOSURE 0.5 0.5 ;

    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 200 ) ( 0.000025 400.00207 ) ( 0.2 416.6 ) ( 0.5 441.5 ) ( 1 483 ) ( 1.5 524.5 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.000025 400.00207 ) ( 0.2 416.6 ) ( 0.5 441.5 ) ( 1 483 ) ( 1.5 524.5 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        TABLEENTRIES	1.666667 ;
    DCCURRENTDENSITY	AVERAGE 1.666667 ; 

END RV

LAYER AP
    TYPE ROUTING ;
    DIRECTION VERTICAL ;
    PITCH   4.500000 4.500000 ;
    OFFSET 0.000000 0.000000 ;
    MINWIDTH	2.000000 ;
    MAXWIDTH	35.000000 ;
    WIDTH   2.000000 ;

    SPACING 2.000000 ;
    HEIGHT  3.105 ;
    THICKNESS	1.450 ;
 
    MINIMUMDENSITY  10 ;
    MAXIMUMDENSITY  70 ;
    DENSITYCHECKWINDOW 100 100 ;
    DENSITYCHECKSTEP	50 ;
 
    ANTENNAMODEL OXIDE1 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 2000 ) ( 0.000025 30000.2 ) ( 0.2 31600.0 ) ( 0.5 34000.0 ) ( 1 38000 ) ( 1.5 42000.0 ) ) ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNADIFFSIDEAREARATIO PWL ( ( 0 1000 ) ( 0.000025 30000.2 ) ( 0.2 31600.0 ) ( 0.5 34000.0 ) ( 1 38000 ) ( 1.5 42000.0 ) ) ;

    
    ACCURRENTDENSITY	AVERAGE
        FREQUENCY	500 ;
        WIDTH    	 1.800000 4.500000 7.200000 13.500000 18.000000 31.500000 ;
        TABLEENTRIES	 3.000000 3.000000 3.000000 3.000000 3.000000 3.000000 ;

    ACCURRENTDENSITY	RMS
        FREQUENCY	500 ;
        WIDTH    	 1.800000 4.500000 7.200000 13.500000 18.000000 31.500000 ;
        TABLEENTRIES	 5.698835 4.539900 4.200498 3.916235 3.831145 3.718884 ;

    ACCURRENTDENSITY	PEAK
        FREQUENCY	500 ;
        WIDTH    	 1.800000 4.500000 7.200000 13.500000 18.000000 31.500000 ;
        TABLEENTRIES	 82.024387 82.024387 82.024387 82.024387 82.024387 82.024387 ;

    DCCURRENTDENSITY	AVERAGE
        WIDTH    	 1.800000 4.500000 7.200000 13.500000 18.000000 31.500000 ;
        TABLEENTRIES	 3.000000 3.000000 3.000000 3.000000 3.000000 3.000000 ;

    RESISTANCE RPERSQ 0.0210000000 ;
    CAPACITANCE CPERSQDIST 0.0000600000 ;
    EDGECAPACITANCE 0.0000591000 ;
END AP

LAYER OVERLAP
	TYPE OVERLAP ;
END OVERLAP

VIA VIA12_square
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
END VIA12_square

VIA VIA12_slot
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.025 0.065 0.025 ;
	LAYER VIA1 ;
		RECT -0.065 -0.025 0.065 0.025 ;
	LAYER M2 ;
		RECT -0.065 -0.025 0.065 0.025 ;
END VIA12_slot

VIA VIA12_slotV
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.065 0.025 0.065 ;
	LAYER VIA1 ;
		RECT -0.025 -0.065 0.025 0.065 ;
	LAYER M2 ;
		RECT -0.025 -0.065 0.025 0.065 ;
END VIA12_slotV

VIA VIA12_1cut DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA12_1cut

VIA VIA12_1cut_FAT_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.075 0.025 0.075 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.075 -0.025 0.075 0.025 ;
END VIA12_1cut_FAT_C

VIA VIA12_1cut_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA12_1cut_H

VIA VIA12_1cut_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA12_1cut_V

VIA VIA12_1cut_EN1415 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA12_1cut_EN1415

VIA VIA12_2cut_P1_CV DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.105 0.025 0.105 ;
	LAYER VIA1 ;
		RECT -0.025 -0.065 0.025 0.065 ;
	LAYER M2 ;
		RECT -0.055 -0.075 0.055 0.075 ;
END VIA12_2cut_P1_CV

VIA VIA12_2cut_P1_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.025 0.155 ;
	LAYER VIA1 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.125 ;
END VIA12_2cut_P1_N

VIA VIA12_2cut_P1_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.155 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M2 ;
		RECT -0.055 -0.125 0.055 0.025 ;
END VIA12_2cut_P1_S

VIA VIA12_2cut_P2_BLC DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.075 -0.055 0.075 0.055 ;
	LAYER VIA1 ;
		RECT -0.065 -0.025 0.065 0.025 ;
	LAYER M2 ;
		RECT -0.22 -0.025 0.22 0.025 ;
END VIA12_2cut_P2_BLC

VIA VIA12_2cut_P2_SLE DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA1 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M2 ;
		RECT -0.065 -0.025 0.375 0.025 ;
END VIA12_2cut_P2_SLE

VIA VIA12_2cut_P2_SLW DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M2 ;
		RECT -0.375 -0.025 0.065 0.025 ;
END VIA12_2cut_P2_SLW

VIA VIA12_2cut_P3_CH DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.075 -0.055 0.075 0.055 ;
	LAYER VIA1 ;
		RECT -0.065 -0.025 0.065 0.025 ;
	LAYER M2 ;
		RECT -0.105 -0.025 0.105 0.025 ;
END VIA12_2cut_P3_CH

VIA VIA12_2cut_P3_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA1 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.155 0.025 ;
END VIA12_2cut_P3_E

VIA VIA12_2cut_P3_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M2 ;
		RECT -0.155 -0.025 0.055 0.025 ;
END VIA12_2cut_P3_W

VIA VIA12_4cut DEFAULT
	RESISTANCE 2.0000000000 ;
	LAYER M1 ;
		RECT -0.09 -0.12 0.09 0.12 ;
	LAYER VIA1 ;
		RECT -0.09 -0.09 -0.04 -0.04 ;
		RECT 0.04 -0.09 0.09 -0.04 ;
		RECT -0.09 0.04 -0.04 0.09 ;
		RECT 0.04 0.04 0.09 0.09 ;
	LAYER M2 ;
		RECT -0.12 -0.09 0.12 0.09 ;
END VIA12_4cut

VIA VIA12_FBD_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.165 0.085 ;
	LAYER VIA1 ;
		RECT 0.005 0.005 0.135 0.055 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.165 0.085 ;
END VIA12_FBD_XEN

VIA VIA12_FBD_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.085 0.165 0.025 ;
	LAYER VIA1 ;
		RECT 0.005 -0.055 0.135 -0.005 ;
	LAYER M2 ;
		RECT -0.025 -0.085 0.165 0.025 ;
END VIA12_FBD_XES

VIA VIA12_FBD_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.165 -0.025 0.025 0.085 ;
	LAYER VIA1 ;
		RECT -0.135 0.005 -0.005 0.055 ;
	LAYER M2 ;
		RECT -0.165 -0.025 0.025 0.085 ;
END VIA12_FBD_XWN

VIA VIA12_FBD_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.165 -0.085 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.135 -0.055 -0.005 -0.005 ;
	LAYER M2 ;
		RECT -0.165 -0.085 0.025 0.025 ;
END VIA12_FBD_XWS

VIA VIA12_FBD_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.085 0.165 ;
	LAYER VIA1 ;
		RECT 0.005 0.005 0.055 0.135 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.085 0.165 ;
END VIA12_FBD_YEN

VIA VIA12_FBD_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.165 0.085 0.025 ;
	LAYER VIA1 ;
		RECT 0.005 -0.135 0.055 -0.005 ;
	LAYER M2 ;
		RECT -0.025 -0.165 0.085 0.025 ;
END VIA12_FBD_YES

VIA VIA12_FBD_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.025 0.025 0.165 ;
	LAYER VIA1 ;
		RECT -0.055 0.005 -0.005 0.135 ;
	LAYER M2 ;
		RECT -0.085 -0.025 0.025 0.165 ;
END VIA12_FBD_YWN

VIA VIA12_FBD_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.165 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.055 -0.135 -0.005 -0.005 ;
	LAYER M2 ;
		RECT -0.085 -0.165 0.025 0.025 ;
END VIA12_FBD_YWS

VIA VIA12_FBS_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.085 0.085 ;
	LAYER VIA1 ;
		RECT 0.005 0.005 0.055 0.055 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.085 0.085 ;
END VIA12_FBS_EN

VIA VIA12_FBS_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.085 0.085 0.025 ;
	LAYER VIA1 ;
		RECT 0.005 -0.055 0.055 -0.005 ;
	LAYER M2 ;
		RECT -0.025 -0.085 0.085 0.025 ;
END VIA12_FBS_ES

VIA VIA12_FBS_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.025 0.025 0.085 ;
	LAYER VIA1 ;
		RECT -0.055 0.005 -0.005 0.055 ;
	LAYER M2 ;
		RECT -0.085 -0.025 0.025 0.085 ;
END VIA12_FBS_WN

VIA VIA12_FBS_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.085 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.055 -0.055 -0.005 -0.005 ;
	LAYER M2 ;
		RECT -0.085 -0.085 0.025 0.025 ;
END VIA12_FBS_WS

VIA VIA12_PBD_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.025 0.175 0.025 ;
	LAYER VIA1 ;
		RECT 0.005 -0.025 0.135 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.055 0.165 0.055 ;
END VIA12_PBD_E

VIA VIA12_PBD_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.035 0.025 0.175 ;
	LAYER VIA1 ;
		RECT -0.025 0.005 0.025 0.135 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.165 ;
END VIA12_PBD_N

VIA VIA12_PBD_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.175 0.025 0.035 ;
	LAYER VIA1 ;
		RECT -0.025 -0.135 0.025 -0.005 ;
	LAYER M2 ;
		RECT -0.055 -0.165 0.055 0.025 ;
END VIA12_PBD_S

VIA VIA12_PBD_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.175 -0.025 0.035 0.025 ;
	LAYER VIA1 ;
		RECT -0.135 -0.025 -0.005 0.025 ;
	LAYER M2 ;
		RECT -0.165 -0.055 0.025 0.055 ;
END VIA12_PBD_W

VIA VIA12_PBS_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA12_PBS_H

VIA VIA12_FBD20_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.145 0.065 ;
	LAYER VIA1 ;
		RECT -0.005 -0.005 0.125 0.045 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.145 0.065 ;
END VIA12_FBD20_XEN

VIA VIA12_FBD20_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.065 0.145 0.025 ;
	LAYER VIA1 ;
		RECT -0.005 -0.045 0.125 0.005 ;
	LAYER M2 ;
		RECT -0.025 -0.065 0.145 0.025 ;
END VIA12_FBD20_XES

VIA VIA12_FBD20_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.145 -0.025 0.025 0.065 ;
	LAYER VIA1 ;
		RECT -0.125 -0.005 0.005 0.045 ;
	LAYER M2 ;
		RECT -0.145 -0.025 0.025 0.065 ;
END VIA12_FBD20_XWN

VIA VIA12_FBD20_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.145 -0.065 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.125 -0.045 0.005 0.005 ;
	LAYER M2 ;
		RECT -0.145 -0.065 0.025 0.025 ;
END VIA12_FBD20_XWS

VIA VIA12_FBD20_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.065 0.145 ;
	LAYER VIA1 ;
		RECT -0.005 -0.005 0.045 0.125 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.065 0.145 ;
END VIA12_FBD20_YEN

VIA VIA12_FBD20_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.145 0.065 0.025 ;
	LAYER VIA1 ;
		RECT -0.005 -0.125 0.045 0.005 ;
	LAYER M2 ;
		RECT -0.025 -0.145 0.065 0.025 ;
END VIA12_FBD20_YES

VIA VIA12_FBD20_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.025 0.025 0.145 ;
	LAYER VIA1 ;
		RECT -0.045 -0.005 0.005 0.125 ;
	LAYER M2 ;
		RECT -0.065 -0.025 0.025 0.145 ;
END VIA12_FBD20_YWN

VIA VIA12_FBD20_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.065 -0.145 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.045 -0.125 0.005 0.005 ;
	LAYER M2 ;
		RECT -0.065 -0.145 0.025 0.025 ;
END VIA12_FBD20_YWS

VIA VIA12_FBD30_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.125 0.085 ;
	LAYER VIA1 ;
		RECT -0.015 0.005 0.115 0.055 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.125 0.085 ;
END VIA12_FBD30_XEN

VIA VIA12_FBD30_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.085 0.125 0.025 ;
	LAYER VIA1 ;
		RECT -0.015 -0.055 0.115 -0.005 ;
	LAYER M2 ;
		RECT -0.025 -0.085 0.125 0.025 ;
END VIA12_FBD30_XES

VIA VIA12_FBD30_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.125 -0.025 0.025 0.085 ;
	LAYER VIA1 ;
		RECT -0.115 0.005 0.015 0.055 ;
	LAYER M2 ;
		RECT -0.125 -0.025 0.025 0.085 ;
END VIA12_FBD30_XWN

VIA VIA12_FBD30_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.125 -0.085 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.115 -0.055 0.015 -0.005 ;
	LAYER M2 ;
		RECT -0.125 -0.085 0.025 0.025 ;
END VIA12_FBD30_XWS

VIA VIA12_FBD30_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.085 0.125 ;
	LAYER VIA1 ;
		RECT 0.005 -0.015 0.055 0.115 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.085 0.125 ;
END VIA12_FBD30_YEN

VIA VIA12_FBD30_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.125 0.085 0.025 ;
	LAYER VIA1 ;
		RECT 0.005 -0.115 0.055 0.015 ;
	LAYER M2 ;
		RECT -0.025 -0.125 0.085 0.025 ;
END VIA12_FBD30_YES

VIA VIA12_FBD30_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.025 0.025 0.125 ;
	LAYER VIA1 ;
		RECT -0.055 -0.015 -0.005 0.115 ;
	LAYER M2 ;
		RECT -0.085 -0.025 0.025 0.125 ;
END VIA12_FBD30_YWN

VIA VIA12_FBD30_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.085 -0.125 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.055 -0.115 -0.005 0.015 ;
	LAYER M2 ;
		RECT -0.085 -0.125 0.025 0.025 ;
END VIA12_FBD30_YWS

VIA VIA12_PBDB_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.005 -0.045 0.165 0.045 ;
	LAYER VIA1 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA12_PBDB_E

VIA VIA12_PBDB_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.045 -0.005 0.045 0.165 ;
	LAYER VIA1 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA12_PBDB_N

VIA VIA12_PBDB_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.045 -0.165 0.045 0.005 ;
	LAYER VIA1 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M2 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA12_PBDB_S

VIA VIA12_PBDB_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.165 -0.045 0.005 0.045 ;
	LAYER VIA1 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M2 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA12_PBDB_W

VIA VIA12_PBDU_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.045 -0.025 0.165 0.025 ;
	LAYER VIA1 ;
		RECT -0.005 -0.025 0.125 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.045 0.145 0.045 ;
END VIA12_PBDU_E

VIA VIA12_PBDU_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.045 0.025 0.165 ;
	LAYER VIA1 ;
		RECT -0.025 -0.005 0.025 0.125 ;
	LAYER M2 ;
		RECT -0.045 -0.025 0.045 0.145 ;
END VIA12_PBDU_N

VIA VIA12_PBDU_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.165 0.025 0.045 ;
	LAYER VIA1 ;
		RECT -0.025 -0.125 0.025 0.005 ;
	LAYER M2 ;
		RECT -0.045 -0.145 0.045 0.025 ;
END VIA12_PBDU_S

VIA VIA12_PBDU_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.165 -0.025 0.045 0.025 ;
	LAYER VIA1 ;
		RECT -0.125 -0.025 0.005 0.025 ;
	LAYER M2 ;
		RECT -0.145 -0.045 0.025 0.045 ;
END VIA12_PBDU_W

VIA VIA12_PBDE_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.185 0.025 ;
	LAYER VIA1 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA12_PBDE_E

VIA VIA12_PBDE_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.025 0.185 ;
	LAYER VIA1 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA12_PBDE_N

VIA VIA12_PBDE_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.185 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M2 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA12_PBDE_S

VIA VIA12_PBDE_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M1 ;
		RECT -0.185 -0.025 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M2 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA12_PBDE_W

VIA VIA12_FBS25_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.025 0.075 0.075 ;
	LAYER VIA1 ;
		RECT 0 0 0.05 0.05 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.075 0.075 ;
END VIA12_FBS25_EN

VIA VIA12_FBS25_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.075 0.075 0.025 ;
	LAYER VIA1 ;
		RECT 0 -0.05 0.05 0 ;
	LAYER M2 ;
		RECT -0.025 -0.075 0.075 0.025 ;
END VIA12_FBS25_ES

VIA VIA12_FBS25_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.075 -0.025 0.025 0.075 ;
	LAYER VIA1 ;
		RECT -0.05 0 0 0.05 ;
	LAYER M2 ;
		RECT -0.075 -0.025 0.025 0.075 ;
END VIA12_FBS25_WN

VIA VIA12_FBS25_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.075 -0.075 0.025 0.025 ;
	LAYER VIA1 ;
		RECT -0.05 -0.05 0 0 ;
	LAYER M2 ;
		RECT -0.075 -0.075 0.025 0.025 ;
END VIA12_FBS25_WS

VIA VIA12_PBSU_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA12_PBSU_H

VIA VIA12_PBSB_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA12_PBSB_H

VIA VIA12_PBS_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA12_PBS_V

VIA VIA12_PBSU_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA12_PBSU_V

VIA VIA12_PBSB_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M1 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA1 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA12_PBSB_V


VIA VIA23_1cut DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA23_1cut

VIA VIA23_1cut_FAT_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.075 -0.025 0.075 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.075 0.025 0.075 ;
END VIA23_1cut_FAT_C

VIA VIA23_1cut_EN1415 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA23_1cut_EN1415

VIA VIA23_1stack_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.14 -0.025 0.14 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA23_1stack_C

VIA VIA23_1stack_E DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.225 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA23_1stack_E

VIA VIA23_1stack_W DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.225 -0.025 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA23_1stack_W

VIA VIA23_2cut_P1_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.155 0.025 ;
	LAYER VIA2 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.125 0.055 ;
END VIA23_2cut_P1_E

VIA VIA23_2cut_P1_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.155 -0.025 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M3 ;
		RECT -0.125 -0.055 0.025 0.055 ;
END VIA23_2cut_P1_W

VIA VIA23_2cut_P2_BLC DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.075 0.055 0.075 ;
	LAYER VIA2 ;
		RECT -0.025 -0.065 0.025 0.065 ;
	LAYER M3 ;
		RECT -0.025 -0.22 0.025 0.22 ;
END VIA23_2cut_P2_BLC

VIA VIA23_2cut_P2_BLN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.125 ;
	LAYER VIA2 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M3 ;
		RECT -0.025 -0.17 0.025 0.27 ;
END VIA23_2cut_P2_BLN

VIA VIA23_2cut_P2_BLS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.125 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M3 ;
		RECT -0.025 -0.27 0.025 0.17 ;
END VIA23_2cut_P2_BLS

VIA VIA23_2cut_P2_SLN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.125 ;
	LAYER VIA2 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M3 ;
		RECT -0.025 -0.065 0.025 0.375 ;
END VIA23_2cut_P2_SLN

VIA VIA23_2cut_P2_SLS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.125 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M3 ;
		RECT -0.025 -0.375 0.025 0.065 ;
END VIA23_2cut_P2_SLS

VIA VIA23_2cut_P3_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.125 ;
	LAYER VIA2 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.155 ;
END VIA23_2cut_P3_N

VIA VIA23_2cut_P3_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.125 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M3 ;
		RECT -0.025 -0.155 0.025 0.055 ;
END VIA23_2cut_P3_S

VIA VIA23_4cut DEFAULT
	RESISTANCE 2.0000000000 ;
	LAYER M2 ;
		RECT -0.12 -0.09 0.12 0.09 ;
	LAYER VIA2 ;
		RECT -0.09 -0.09 -0.04 -0.04 ;
		RECT 0.04 -0.09 0.09 -0.04 ;
		RECT -0.09 0.04 -0.04 0.09 ;
		RECT 0.04 0.04 0.09 0.09 ;
	LAYER M3 ;
		RECT -0.09 -0.12 0.09 0.12 ;
END VIA23_4cut

VIA VIA23_FBD_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.165 0.085 ;
	LAYER VIA2 ;
		RECT 0.005 0.005 0.135 0.055 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.165 0.085 ;
END VIA23_FBD_XEN

VIA VIA23_FBD_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.085 0.165 0.025 ;
	LAYER VIA2 ;
		RECT 0.005 -0.055 0.135 -0.005 ;
	LAYER M3 ;
		RECT -0.025 -0.085 0.165 0.025 ;
END VIA23_FBD_XES

VIA VIA23_FBD_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.165 -0.025 0.025 0.085 ;
	LAYER VIA2 ;
		RECT -0.135 0.005 -0.005 0.055 ;
	LAYER M3 ;
		RECT -0.165 -0.025 0.025 0.085 ;
END VIA23_FBD_XWN

VIA VIA23_FBD_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.165 -0.085 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.135 -0.055 -0.005 -0.005 ;
	LAYER M3 ;
		RECT -0.165 -0.085 0.025 0.025 ;
END VIA23_FBD_XWS

VIA VIA23_FBD_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.085 0.165 ;
	LAYER VIA2 ;
		RECT 0.005 0.005 0.055 0.135 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.085 0.165 ;
END VIA23_FBD_YEN

VIA VIA23_FBD_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.165 0.085 0.025 ;
	LAYER VIA2 ;
		RECT 0.005 -0.135 0.055 -0.005 ;
	LAYER M3 ;
		RECT -0.025 -0.165 0.085 0.025 ;
END VIA23_FBD_YES

VIA VIA23_FBD_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.085 -0.025 0.025 0.165 ;
	LAYER VIA2 ;
		RECT -0.055 0.005 -0.005 0.135 ;
	LAYER M3 ;
		RECT -0.085 -0.025 0.025 0.165 ;
END VIA23_FBD_YWN

VIA VIA23_FBD_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.085 -0.165 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.055 -0.135 -0.005 -0.005 ;
	LAYER M3 ;
		RECT -0.085 -0.165 0.025 0.025 ;
END VIA23_FBD_YWS

VIA VIA23_FBS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.055 0.055 0.055 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA23_FBS

VIA VIA23_FBS_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.085 0.085 ;
	LAYER VIA2 ;
		RECT 0.005 0.005 0.055 0.055 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.085 0.085 ;
END VIA23_FBS_EN

VIA VIA23_FBS_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.085 0.085 0.025 ;
	LAYER VIA2 ;
		RECT 0.005 -0.055 0.055 -0.005 ;
	LAYER M3 ;
		RECT -0.025 -0.085 0.085 0.025 ;
END VIA23_FBS_ES

VIA VIA23_FBS_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.085 -0.025 0.025 0.085 ;
	LAYER VIA2 ;
		RECT -0.055 0.005 -0.005 0.055 ;
	LAYER M3 ;
		RECT -0.085 -0.025 0.025 0.085 ;
END VIA23_FBS_WN

VIA VIA23_FBS_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.085 -0.085 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.055 -0.055 -0.005 -0.005 ;
	LAYER M3 ;
		RECT -0.085 -0.085 0.025 0.025 ;
END VIA23_FBS_WS

VIA VIA23_PBD_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.025 0.175 0.025 ;
	LAYER VIA2 ;
		RECT 0.005 -0.025 0.135 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.165 0.055 ;
END VIA23_PBD_E

VIA VIA23_PBD_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.035 0.025 0.175 ;
	LAYER VIA2 ;
		RECT -0.025 0.005 0.025 0.135 ;
	LAYER M3 ;
		RECT -0.055 -0.025 0.055 0.165 ;
END VIA23_PBD_N

VIA VIA23_PBD_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.175 0.025 0.035 ;
	LAYER VIA2 ;
		RECT -0.025 -0.135 0.025 -0.005 ;
	LAYER M3 ;
		RECT -0.055 -0.165 0.055 0.025 ;
END VIA23_PBD_S

VIA VIA23_PBD_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.175 -0.025 0.035 0.025 ;
	LAYER VIA2 ;
		RECT -0.135 -0.025 -0.005 0.025 ;
	LAYER M3 ;
		RECT -0.165 -0.055 0.025 0.055 ;
END VIA23_PBD_W

VIA VIA23_PBS_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA23_PBS_H

VIA VIA23_PBS_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA23_PBS_V

VIA VIA23_FBD20_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.145 0.065 ;
	LAYER VIA2 ;
		RECT -0.005 -0.005 0.125 0.045 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.145 0.065 ;
END VIA23_FBD20_XEN

VIA VIA23_FBD20_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.065 0.145 0.025 ;
	LAYER VIA2 ;
		RECT -0.005 -0.045 0.125 0.005 ;
	LAYER M3 ;
		RECT -0.025 -0.065 0.145 0.025 ;
END VIA23_FBD20_XES

VIA VIA23_FBD20_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.145 -0.025 0.025 0.065 ;
	LAYER VIA2 ;
		RECT -0.125 -0.005 0.005 0.045 ;
	LAYER M3 ;
		RECT -0.145 -0.025 0.025 0.065 ;
END VIA23_FBD20_XWN

VIA VIA23_FBD20_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.145 -0.065 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.125 -0.045 0.005 0.005 ;
	LAYER M3 ;
		RECT -0.145 -0.065 0.025 0.025 ;
END VIA23_FBD20_XWS

VIA VIA23_FBD20_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.065 0.145 ;
	LAYER VIA2 ;
		RECT -0.005 -0.005 0.045 0.125 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.065 0.145 ;
END VIA23_FBD20_YEN

VIA VIA23_FBD20_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.145 0.065 0.025 ;
	LAYER VIA2 ;
		RECT -0.005 -0.125 0.045 0.005 ;
	LAYER M3 ;
		RECT -0.025 -0.145 0.065 0.025 ;
END VIA23_FBD20_YES

VIA VIA23_FBD20_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.065 -0.025 0.025 0.145 ;
	LAYER VIA2 ;
		RECT -0.045 -0.005 0.005 0.125 ;
	LAYER M3 ;
		RECT -0.065 -0.025 0.025 0.145 ;
END VIA23_FBD20_YWN

VIA VIA23_FBD20_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.065 -0.145 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.045 -0.125 0.005 0.005 ;
	LAYER M3 ;
		RECT -0.065 -0.145 0.025 0.025 ;
END VIA23_FBD20_YWS

VIA VIA23_FBD30_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.125 0.085 ;
	LAYER VIA2 ;
		RECT -0.015 0.005 0.115 0.055 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.125 0.085 ;
END VIA23_FBD30_XEN

VIA VIA23_FBD30_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.085 0.125 0.025 ;
	LAYER VIA2 ;
		RECT -0.015 -0.055 0.115 -0.005 ;
	LAYER M3 ;
		RECT -0.025 -0.085 0.125 0.025 ;
END VIA23_FBD30_XES

VIA VIA23_FBD30_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.125 -0.025 0.025 0.085 ;
	LAYER VIA2 ;
		RECT -0.115 0.005 0.015 0.055 ;
	LAYER M3 ;
		RECT -0.125 -0.025 0.025 0.085 ;
END VIA23_FBD30_XWN

VIA VIA23_FBD30_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.125 -0.085 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.115 -0.055 0.015 -0.005 ;
	LAYER M3 ;
		RECT -0.125 -0.085 0.025 0.025 ;
END VIA23_FBD30_XWS

VIA VIA23_FBD30_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.085 0.125 ;
	LAYER VIA2 ;
		RECT 0.005 -0.015 0.055 0.115 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.085 0.125 ;
END VIA23_FBD30_YEN

VIA VIA23_FBD30_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.125 0.085 0.025 ;
	LAYER VIA2 ;
		RECT 0.005 -0.115 0.055 0.015 ;
	LAYER M3 ;
		RECT -0.025 -0.125 0.085 0.025 ;
END VIA23_FBD30_YES

VIA VIA23_FBD30_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.085 -0.025 0.025 0.125 ;
	LAYER VIA2 ;
		RECT -0.055 -0.015 -0.005 0.115 ;
	LAYER M3 ;
		RECT -0.085 -0.025 0.025 0.125 ;
END VIA23_FBD30_YWN

VIA VIA23_FBD30_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.085 -0.125 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.055 -0.115 -0.005 0.015 ;
	LAYER M3 ;
		RECT -0.085 -0.125 0.025 0.025 ;
END VIA23_FBD30_YWS

VIA VIA23_PBDB_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.005 -0.045 0.165 0.045 ;
	LAYER VIA2 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA23_PBDB_E

VIA VIA23_PBDB_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.045 -0.005 0.045 0.165 ;
	LAYER VIA2 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA23_PBDB_N

VIA VIA23_PBDB_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.045 -0.165 0.045 0.005 ;
	LAYER VIA2 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M3 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA23_PBDB_S

VIA VIA23_PBDB_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.165 -0.045 0.005 0.045 ;
	LAYER VIA2 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M3 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA23_PBDB_W

VIA VIA23_PBDU_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.045 -0.025 0.165 0.025 ;
	LAYER VIA2 ;
		RECT -0.005 -0.025 0.125 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.045 0.145 0.045 ;
END VIA23_PBDU_E

VIA VIA23_PBDU_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.045 0.025 0.165 ;
	LAYER VIA2 ;
		RECT -0.025 -0.005 0.025 0.125 ;
	LAYER M3 ;
		RECT -0.045 -0.025 0.045 0.145 ;
END VIA23_PBDU_N

VIA VIA23_PBDU_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.165 0.025 0.045 ;
	LAYER VIA2 ;
		RECT -0.025 -0.125 0.025 0.005 ;
	LAYER M3 ;
		RECT -0.045 -0.145 0.045 0.025 ;
END VIA23_PBDU_S

VIA VIA23_PBDU_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.165 -0.025 0.045 0.025 ;
	LAYER VIA2 ;
		RECT -0.125 -0.025 0.005 0.025 ;
	LAYER M3 ;
		RECT -0.145 -0.045 0.025 0.045 ;
END VIA23_PBDU_W

VIA VIA23_PBDE_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.185 0.025 ;
	LAYER VIA2 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA23_PBDE_E

VIA VIA23_PBDE_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.025 0.185 ;
	LAYER VIA2 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA23_PBDE_N

VIA VIA23_PBDE_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.185 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M3 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA23_PBDE_S

VIA VIA23_PBDE_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M2 ;
		RECT -0.185 -0.025 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M3 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA23_PBDE_W

VIA VIA23_FBS25 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.05 -0.05 0.05 0.05 ;
END VIA23_FBS25

VIA VIA23_FBS25_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.025 0.075 0.075 ;
	LAYER VIA2 ;
		RECT 0 0 0.05 0.05 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.075 0.075 ;
END VIA23_FBS25_EN

VIA VIA23_FBS25_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.075 0.075 0.025 ;
	LAYER VIA2 ;
		RECT 0 -0.05 0.05 0 ;
	LAYER M3 ;
		RECT -0.025 -0.075 0.075 0.025 ;
END VIA23_FBS25_ES

VIA VIA23_FBS25_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.075 -0.025 0.025 0.075 ;
	LAYER VIA2 ;
		RECT -0.05 0 0 0.05 ;
	LAYER M3 ;
		RECT -0.075 -0.025 0.025 0.075 ;
END VIA23_FBS25_WN

VIA VIA23_FBS25_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.075 -0.075 0.025 0.025 ;
	LAYER VIA2 ;
		RECT -0.05 -0.05 0 0 ;
	LAYER M3 ;
		RECT -0.075 -0.075 0.025 0.025 ;
END VIA23_FBS25_WS

VIA VIA23_PBSU_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA23_PBSU_H

VIA VIA23_PBSU_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA23_PBSU_V

VIA VIA23_PBSB_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA23_PBSB_H

VIA VIA23_PBSB_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M2 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA2 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M3 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA23_PBSB_V


VIA VIA34_1cut DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA34_1cut

VIA VIA34_1cut_FAT_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.075 0.025 0.075 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.075 -0.025 0.075 0.025 ;
END VIA34_1cut_FAT_C

VIA VIA34_1cut_EN1415 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA34_1cut_EN1415

VIA VIA34_1stack_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.17 0.025 0.17 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA34_1stack_C

VIA VIA34_1stack_N DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.285 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA34_1stack_N

VIA VIA34_1stack_S DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.285 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA34_1stack_S

VIA VIA34_2cut_P1_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.155 ;
	LAYER VIA3 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.125 ;
END VIA34_2cut_P1_N

VIA VIA34_2cut_P1_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.155 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M4 ;
		RECT -0.055 -0.125 0.055 0.025 ;
END VIA34_2cut_P1_S

VIA VIA34_2cut_P2_BLC DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.075 -0.055 0.075 0.055 ;
	LAYER VIA3 ;
		RECT -0.065 -0.025 0.065 0.025 ;
	LAYER M4 ;
		RECT -0.22 -0.025 0.22 0.025 ;
END VIA34_2cut_P2_BLC

VIA VIA34_2cut_P2_BLE DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA3 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M4 ;
		RECT -0.17 -0.025 0.27 0.025 ;
END VIA34_2cut_P2_BLE

VIA VIA34_2cut_P2_BLW DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M4 ;
		RECT -0.27 -0.025 0.17 0.025 ;
END VIA34_2cut_P2_BLW

VIA VIA34_2cut_P2_SLE DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA3 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M4 ;
		RECT -0.065 -0.025 0.375 0.025 ;
END VIA34_2cut_P2_SLE

VIA VIA34_2cut_P2_SLW DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M4 ;
		RECT -0.375 -0.025 0.065 0.025 ;
END VIA34_2cut_P2_SLW

VIA VIA34_2cut_P3_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA3 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.155 0.025 ;
END VIA34_2cut_P3_E

VIA VIA34_2cut_P3_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M4 ;
		RECT -0.155 -0.025 0.055 0.025 ;
END VIA34_2cut_P3_W

VIA VIA34_4cut DEFAULT
	RESISTANCE 2.0000000000 ;
	LAYER M3 ;
		RECT -0.09 -0.12 0.09 0.12 ;
	LAYER VIA3 ;
		RECT -0.09 -0.09 -0.04 -0.04 ;
		RECT 0.04 -0.09 0.09 -0.04 ;
		RECT -0.09 0.04 -0.04 0.09 ;
		RECT 0.04 0.04 0.09 0.09 ;
	LAYER M4 ;
		RECT -0.12 -0.09 0.12 0.09 ;
END VIA34_4cut

VIA VIA34_FBD_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.165 0.085 ;
	LAYER VIA3 ;
		RECT 0.005 0.005 0.135 0.055 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.165 0.085 ;
END VIA34_FBD_XEN

VIA VIA34_FBD_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.085 0.165 0.025 ;
	LAYER VIA3 ;
		RECT 0.005 -0.055 0.135 -0.005 ;
	LAYER M4 ;
		RECT -0.025 -0.085 0.165 0.025 ;
END VIA34_FBD_XES

VIA VIA34_FBD_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.165 -0.025 0.025 0.085 ;
	LAYER VIA3 ;
		RECT -0.135 0.005 -0.005 0.055 ;
	LAYER M4 ;
		RECT -0.165 -0.025 0.025 0.085 ;
END VIA34_FBD_XWN

VIA VIA34_FBD_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.165 -0.085 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.135 -0.055 -0.005 -0.005 ;
	LAYER M4 ;
		RECT -0.165 -0.085 0.025 0.025 ;
END VIA34_FBD_XWS

VIA VIA34_FBD_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.085 0.165 ;
	LAYER VIA3 ;
		RECT 0.005 0.005 0.055 0.135 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.085 0.165 ;
END VIA34_FBD_YEN

VIA VIA34_FBD_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.165 0.085 0.025 ;
	LAYER VIA3 ;
		RECT 0.005 -0.135 0.055 -0.005 ;
	LAYER M4 ;
		RECT -0.025 -0.165 0.085 0.025 ;
END VIA34_FBD_YES

VIA VIA34_FBD_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.025 0.025 0.165 ;
	LAYER VIA3 ;
		RECT -0.055 0.005 -0.005 0.135 ;
	LAYER M4 ;
		RECT -0.085 -0.025 0.025 0.165 ;
END VIA34_FBD_YWN

VIA VIA34_FBD_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.165 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.055 -0.135 -0.005 -0.005 ;
	LAYER M4 ;
		RECT -0.085 -0.165 0.025 0.025 ;
END VIA34_FBD_YWS

VIA VIA34_FBS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.055 -0.055 0.055 0.055 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA34_FBS

VIA VIA34_FBS_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.085 0.085 ;
	LAYER VIA3 ;
		RECT 0.005 0.005 0.055 0.055 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.085 0.085 ;
END VIA34_FBS_EN

VIA VIA34_FBS_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.085 0.085 0.025 ;
	LAYER VIA3 ;
		RECT 0.005 -0.055 0.055 -0.005 ;
	LAYER M4 ;
		RECT -0.025 -0.085 0.085 0.025 ;
END VIA34_FBS_ES

VIA VIA34_FBS_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.025 0.025 0.085 ;
	LAYER VIA3 ;
		RECT -0.055 0.005 -0.005 0.055 ;
	LAYER M4 ;
		RECT -0.085 -0.025 0.025 0.085 ;
END VIA34_FBS_WN

VIA VIA34_FBS_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.085 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.055 -0.055 -0.005 -0.005 ;
	LAYER M4 ;
		RECT -0.085 -0.085 0.025 0.025 ;
END VIA34_FBS_WS

VIA VIA34_PBD_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.035 -0.025 0.175 0.025 ;
	LAYER VIA3 ;
		RECT 0.005 -0.025 0.135 0.025 ;
	LAYER M4 ;
		RECT -0.025 -0.055 0.165 0.055 ;
END VIA34_PBD_E

VIA VIA34_PBD_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.035 0.025 0.175 ;
	LAYER VIA3 ;
		RECT -0.025 0.005 0.025 0.135 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.165 ;
END VIA34_PBD_N

VIA VIA34_PBD_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.175 0.025 0.035 ;
	LAYER VIA3 ;
		RECT -0.025 -0.135 0.025 -0.005 ;
	LAYER M4 ;
		RECT -0.055 -0.165 0.055 0.025 ;
END VIA34_PBD_S

VIA VIA34_PBD_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.175 -0.025 0.035 0.025 ;
	LAYER VIA3 ;
		RECT -0.135 -0.025 -0.005 0.025 ;
	LAYER M4 ;
		RECT -0.165 -0.055 0.025 0.055 ;
END VIA34_PBD_W

VIA VIA34_PBS_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA34_PBS_H

VIA VIA34_PBS_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA34_PBS_V

VIA VIA34_FBD20_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.145 0.065 ;
	LAYER VIA3 ;
		RECT -0.005 -0.005 0.125 0.045 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.145 0.065 ;
END VIA34_FBD20_XEN

VIA VIA34_FBD20_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.065 0.145 0.025 ;
	LAYER VIA3 ;
		RECT -0.005 -0.045 0.125 0.005 ;
	LAYER M4 ;
		RECT -0.025 -0.065 0.145 0.025 ;
END VIA34_FBD20_XES

VIA VIA34_FBD20_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.145 -0.025 0.025 0.065 ;
	LAYER VIA3 ;
		RECT -0.125 -0.005 0.005 0.045 ;
	LAYER M4 ;
		RECT -0.145 -0.025 0.025 0.065 ;
END VIA34_FBD20_XWN

VIA VIA34_FBD20_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.145 -0.065 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.125 -0.045 0.005 0.005 ;
	LAYER M4 ;
		RECT -0.145 -0.065 0.025 0.025 ;
END VIA34_FBD20_XWS

VIA VIA34_FBD20_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.065 0.145 ;
	LAYER VIA3 ;
		RECT -0.005 -0.005 0.045 0.125 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.065 0.145 ;
END VIA34_FBD20_YEN

VIA VIA34_FBD20_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.145 0.065 0.025 ;
	LAYER VIA3 ;
		RECT -0.005 -0.125 0.045 0.005 ;
	LAYER M4 ;
		RECT -0.025 -0.145 0.065 0.025 ;
END VIA34_FBD20_YES

VIA VIA34_FBD20_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.065 -0.025 0.025 0.145 ;
	LAYER VIA3 ;
		RECT -0.045 -0.005 0.005 0.125 ;
	LAYER M4 ;
		RECT -0.065 -0.025 0.025 0.145 ;
END VIA34_FBD20_YWN

VIA VIA34_FBD20_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.065 -0.145 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.045 -0.125 0.005 0.005 ;
	LAYER M4 ;
		RECT -0.065 -0.145 0.025 0.025 ;
END VIA34_FBD20_YWS

VIA VIA34_FBD30_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.125 0.085 ;
	LAYER VIA3 ;
		RECT -0.015 0.005 0.115 0.055 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.125 0.085 ;
END VIA34_FBD30_XEN

VIA VIA34_FBD30_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.085 0.125 0.025 ;
	LAYER VIA3 ;
		RECT -0.015 -0.055 0.115 -0.005 ;
	LAYER M4 ;
		RECT -0.025 -0.085 0.125 0.025 ;
END VIA34_FBD30_XES

VIA VIA34_FBD30_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.125 -0.025 0.025 0.085 ;
	LAYER VIA3 ;
		RECT -0.115 0.005 0.015 0.055 ;
	LAYER M4 ;
		RECT -0.125 -0.025 0.025 0.085 ;
END VIA34_FBD30_XWN

VIA VIA34_FBD30_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.125 -0.085 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.115 -0.055 0.015 -0.005 ;
	LAYER M4 ;
		RECT -0.125 -0.085 0.025 0.025 ;
END VIA34_FBD30_XWS

VIA VIA34_FBD30_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.085 0.125 ;
	LAYER VIA3 ;
		RECT 0.005 -0.015 0.055 0.115 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.085 0.125 ;
END VIA34_FBD30_YEN

VIA VIA34_FBD30_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.125 0.085 0.025 ;
	LAYER VIA3 ;
		RECT 0.005 -0.115 0.055 0.015 ;
	LAYER M4 ;
		RECT -0.025 -0.125 0.085 0.025 ;
END VIA34_FBD30_YES

VIA VIA34_FBD30_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.025 0.025 0.125 ;
	LAYER VIA3 ;
		RECT -0.055 -0.015 -0.005 0.115 ;
	LAYER M4 ;
		RECT -0.085 -0.025 0.025 0.125 ;
END VIA34_FBD30_YWN

VIA VIA34_FBD30_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.085 -0.125 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.055 -0.115 -0.005 0.015 ;
	LAYER M4 ;
		RECT -0.085 -0.125 0.025 0.025 ;
END VIA34_FBD30_YWS

VIA VIA34_PBDB_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.005 -0.045 0.165 0.045 ;
	LAYER VIA3 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA34_PBDB_E

VIA VIA34_PBDB_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.045 -0.005 0.045 0.165 ;
	LAYER VIA3 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA34_PBDB_N

VIA VIA34_PBDB_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.045 -0.165 0.045 0.005 ;
	LAYER VIA3 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M4 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA34_PBDB_S

VIA VIA34_PBDB_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.165 -0.045 0.005 0.045 ;
	LAYER VIA3 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M4 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA34_PBDB_W

VIA VIA34_PBDU_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.045 -0.025 0.165 0.025 ;
	LAYER VIA3 ;
		RECT -0.005 -0.025 0.125 0.025 ;
	LAYER M4 ;
		RECT -0.025 -0.045 0.145 0.045 ;
END VIA34_PBDU_E

VIA VIA34_PBDU_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.045 0.025 0.165 ;
	LAYER VIA3 ;
		RECT -0.025 -0.005 0.025 0.125 ;
	LAYER M4 ;
		RECT -0.045 -0.025 0.045 0.145 ;
END VIA34_PBDU_N

VIA VIA34_PBDU_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.165 0.025 0.045 ;
	LAYER VIA3 ;
		RECT -0.025 -0.125 0.025 0.005 ;
	LAYER M4 ;
		RECT -0.045 -0.145 0.045 0.025 ;
END VIA34_PBDU_S

VIA VIA34_PBDU_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.165 -0.025 0.045 0.025 ;
	LAYER VIA3 ;
		RECT -0.125 -0.025 0.005 0.025 ;
	LAYER M4 ;
		RECT -0.145 -0.045 0.025 0.045 ;
END VIA34_PBDU_W

VIA VIA34_PBDE_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.185 0.025 ;
	LAYER VIA3 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA34_PBDE_E

VIA VIA34_PBDE_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.025 0.185 ;
	LAYER VIA3 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA34_PBDE_N

VIA VIA34_PBDE_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.185 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M4 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA34_PBDE_S

VIA VIA34_PBDE_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M3 ;
		RECT -0.185 -0.025 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M4 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA34_PBDE_W

VIA VIA34_FBS25 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.05 -0.05 0.05 0.05 ;
END VIA34_FBS25

VIA VIA34_FBS25_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.025 0.075 0.075 ;
	LAYER VIA3 ;
		RECT 0 0 0.05 0.05 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.075 0.075 ;
END VIA34_FBS25_EN

VIA VIA34_FBS25_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.075 0.075 0.025 ;
	LAYER VIA3 ;
		RECT 0 -0.05 0.05 0 ;
	LAYER M4 ;
		RECT -0.025 -0.075 0.075 0.025 ;
END VIA34_FBS25_ES

VIA VIA34_FBS25_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.075 -0.025 0.025 0.075 ;
	LAYER VIA3 ;
		RECT -0.05 0 0 0.05 ;
	LAYER M4 ;
		RECT -0.075 -0.025 0.025 0.075 ;
END VIA34_FBS25_WN

VIA VIA34_FBS25_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.075 -0.075 0.025 0.025 ;
	LAYER VIA3 ;
		RECT -0.05 -0.05 0 0 ;
	LAYER M4 ;
		RECT -0.075 -0.075 0.025 0.025 ;
END VIA34_FBS25_WS

VIA VIA34_PBSU_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA34_PBSU_H

VIA VIA34_PBSU_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA34_PBSU_V

VIA VIA34_PBSB_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA34_PBSB_H

VIA VIA34_PBSB_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M3 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA3 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA34_PBSB_V


VIA VIA45_1cut DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA45_1cut

VIA VIA45_1cut_FAT_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.075 -0.025 0.075 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.075 0.025 0.075 ;
END VIA45_1cut_FAT_C

VIA VIA45_1cut_EN1415 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA45_1cut_EN1415

VIA VIA45_1stack_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.17 -0.025 0.17 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA45_1stack_C

VIA VIA45_1stack_E DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.285 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA45_1stack_E

VIA VIA45_1stack_W DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.285 -0.025 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA45_1stack_W

VIA VIA45_2cut_P1_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.155 0.025 ;
	LAYER VIA4 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.125 0.055 ;
END VIA45_2cut_P1_E

VIA VIA45_2cut_P1_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.155 -0.025 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M5 ;
		RECT -0.125 -0.055 0.025 0.055 ;
END VIA45_2cut_P1_W

VIA VIA45_2cut_P2_BLC DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.075 0.055 0.075 ;
	LAYER VIA4 ;
		RECT -0.025 -0.065 0.025 0.065 ;
	LAYER M5 ;
		RECT -0.025 -0.22 0.025 0.22 ;
END VIA45_2cut_P2_BLC

VIA VIA45_2cut_P2_BLN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.125 ;
	LAYER VIA4 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M5 ;
		RECT -0.025 -0.17 0.025 0.27 ;
END VIA45_2cut_P2_BLN

VIA VIA45_2cut_P2_BLS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.125 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M5 ;
		RECT -0.025 -0.27 0.025 0.17 ;
END VIA45_2cut_P2_BLS

VIA VIA45_2cut_P2_SLN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.125 ;
	LAYER VIA4 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M5 ;
		RECT -0.025 -0.065 0.025 0.375 ;
END VIA45_2cut_P2_SLN

VIA VIA45_2cut_P2_SLS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.125 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M5 ;
		RECT -0.025 -0.375 0.025 0.065 ;
END VIA45_2cut_P2_SLS

VIA VIA45_2cut_P3_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.125 ;
	LAYER VIA4 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.155 ;
END VIA45_2cut_P3_N

VIA VIA45_2cut_P3_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.125 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M5 ;
		RECT -0.025 -0.155 0.025 0.055 ;
END VIA45_2cut_P3_S

VIA VIA45_4cut DEFAULT
	RESISTANCE 2.0000000000 ;
	LAYER M4 ;
		RECT -0.12 -0.09 0.12 0.09 ;
	LAYER VIA4 ;
		RECT -0.09 -0.09 -0.04 -0.04 ;
		RECT 0.04 -0.09 0.09 -0.04 ;
		RECT -0.09 0.04 -0.04 0.09 ;
		RECT 0.04 0.04 0.09 0.09 ;
	LAYER M5 ;
		RECT -0.09 -0.12 0.09 0.12 ;
END VIA45_4cut

VIA VIA45_FBD_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.165 0.085 ;
	LAYER VIA4 ;
		RECT 0.005 0.005 0.135 0.055 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.165 0.085 ;
END VIA45_FBD_XEN

VIA VIA45_FBD_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.085 0.165 0.025 ;
	LAYER VIA4 ;
		RECT 0.005 -0.055 0.135 -0.005 ;
	LAYER M5 ;
		RECT -0.025 -0.085 0.165 0.025 ;
END VIA45_FBD_XES

VIA VIA45_FBD_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.165 -0.025 0.025 0.085 ;
	LAYER VIA4 ;
		RECT -0.135 0.005 -0.005 0.055 ;
	LAYER M5 ;
		RECT -0.165 -0.025 0.025 0.085 ;
END VIA45_FBD_XWN

VIA VIA45_FBD_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.165 -0.085 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.135 -0.055 -0.005 -0.005 ;
	LAYER M5 ;
		RECT -0.165 -0.085 0.025 0.025 ;
END VIA45_FBD_XWS

VIA VIA45_FBD_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.085 0.165 ;
	LAYER VIA4 ;
		RECT 0.005 0.005 0.055 0.135 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.085 0.165 ;
END VIA45_FBD_YEN

VIA VIA45_FBD_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.165 0.085 0.025 ;
	LAYER VIA4 ;
		RECT 0.005 -0.135 0.055 -0.005 ;
	LAYER M5 ;
		RECT -0.025 -0.165 0.085 0.025 ;
END VIA45_FBD_YES

VIA VIA45_FBD_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.085 -0.025 0.025 0.165 ;
	LAYER VIA4 ;
		RECT -0.055 0.005 -0.005 0.135 ;
	LAYER M5 ;
		RECT -0.085 -0.025 0.025 0.165 ;
END VIA45_FBD_YWN

VIA VIA45_FBD_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.085 -0.165 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.055 -0.135 -0.005 -0.005 ;
	LAYER M5 ;
		RECT -0.085 -0.165 0.025 0.025 ;
END VIA45_FBD_YWS

VIA VIA45_FBS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.055 0.055 0.055 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA45_FBS

VIA VIA45_FBS_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.085 0.085 ;
	LAYER VIA4 ;
		RECT 0.005 0.005 0.055 0.055 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.085 0.085 ;
END VIA45_FBS_EN

VIA VIA45_FBS_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.085 0.085 0.025 ;
	LAYER VIA4 ;
		RECT 0.005 -0.055 0.055 -0.005 ;
	LAYER M5 ;
		RECT -0.025 -0.085 0.085 0.025 ;
END VIA45_FBS_ES

VIA VIA45_FBS_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.085 -0.025 0.025 0.085 ;
	LAYER VIA4 ;
		RECT -0.055 0.005 -0.005 0.055 ;
	LAYER M5 ;
		RECT -0.085 -0.025 0.025 0.085 ;
END VIA45_FBS_WN

VIA VIA45_FBS_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.085 -0.085 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.055 -0.055 -0.005 -0.005 ;
	LAYER M5 ;
		RECT -0.085 -0.085 0.025 0.025 ;
END VIA45_FBS_WS

VIA VIA45_PBD_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.025 0.175 0.025 ;
	LAYER VIA4 ;
		RECT 0.005 -0.025 0.135 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.165 0.055 ;
END VIA45_PBD_E

VIA VIA45_PBD_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.035 0.025 0.175 ;
	LAYER VIA4 ;
		RECT -0.025 0.005 0.025 0.135 ;
	LAYER M5 ;
		RECT -0.055 -0.025 0.055 0.165 ;
END VIA45_PBD_N

VIA VIA45_PBD_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.175 0.025 0.035 ;
	LAYER VIA4 ;
		RECT -0.025 -0.135 0.025 -0.005 ;
	LAYER M5 ;
		RECT -0.055 -0.165 0.055 0.025 ;
END VIA45_PBD_S

VIA VIA45_PBD_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.175 -0.025 0.035 0.025 ;
	LAYER VIA4 ;
		RECT -0.135 -0.025 -0.005 0.025 ;
	LAYER M5 ;
		RECT -0.165 -0.055 0.025 0.055 ;
END VIA45_PBD_W

VIA VIA45_PBS_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA45_PBS_H

VIA VIA45_PBS_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA45_PBS_V

VIA VIA45_FBD20_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.145 0.065 ;
	LAYER VIA4 ;
		RECT -0.005 -0.005 0.125 0.045 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.145 0.065 ;
END VIA45_FBD20_XEN

VIA VIA45_FBD20_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.065 0.145 0.025 ;
	LAYER VIA4 ;
		RECT -0.005 -0.045 0.125 0.005 ;
	LAYER M5 ;
		RECT -0.025 -0.065 0.145 0.025 ;
END VIA45_FBD20_XES

VIA VIA45_FBD20_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.145 -0.025 0.025 0.065 ;
	LAYER VIA4 ;
		RECT -0.125 -0.005 0.005 0.045 ;
	LAYER M5 ;
		RECT -0.145 -0.025 0.025 0.065 ;
END VIA45_FBD20_XWN

VIA VIA45_FBD20_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.145 -0.065 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.125 -0.045 0.005 0.005 ;
	LAYER M5 ;
		RECT -0.145 -0.065 0.025 0.025 ;
END VIA45_FBD20_XWS

VIA VIA45_FBD20_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.065 0.145 ;
	LAYER VIA4 ;
		RECT -0.005 -0.005 0.045 0.125 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.065 0.145 ;
END VIA45_FBD20_YEN

VIA VIA45_FBD20_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.145 0.065 0.025 ;
	LAYER VIA4 ;
		RECT -0.005 -0.125 0.045 0.005 ;
	LAYER M5 ;
		RECT -0.025 -0.145 0.065 0.025 ;
END VIA45_FBD20_YES

VIA VIA45_FBD20_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.065 -0.025 0.025 0.145 ;
	LAYER VIA4 ;
		RECT -0.045 -0.005 0.005 0.125 ;
	LAYER M5 ;
		RECT -0.065 -0.025 0.025 0.145 ;
END VIA45_FBD20_YWN

VIA VIA45_FBD20_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.065 -0.145 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.045 -0.125 0.005 0.005 ;
	LAYER M5 ;
		RECT -0.065 -0.145 0.025 0.025 ;
END VIA45_FBD20_YWS

VIA VIA45_FBD30_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.125 0.085 ;
	LAYER VIA4 ;
		RECT -0.015 0.005 0.115 0.055 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.125 0.085 ;
END VIA45_FBD30_XEN

VIA VIA45_FBD30_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.085 0.125 0.025 ;
	LAYER VIA4 ;
		RECT -0.015 -0.055 0.115 -0.005 ;
	LAYER M5 ;
		RECT -0.025 -0.085 0.125 0.025 ;
END VIA45_FBD30_XES

VIA VIA45_FBD30_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.125 -0.025 0.025 0.085 ;
	LAYER VIA4 ;
		RECT -0.115 0.005 0.015 0.055 ;
	LAYER M5 ;
		RECT -0.125 -0.025 0.025 0.085 ;
END VIA45_FBD30_XWN

VIA VIA45_FBD30_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.125 -0.085 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.115 -0.055 0.015 -0.005 ;
	LAYER M5 ;
		RECT -0.125 -0.085 0.025 0.025 ;
END VIA45_FBD30_XWS

VIA VIA45_FBD30_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.085 0.125 ;
	LAYER VIA4 ;
		RECT 0.005 -0.015 0.055 0.115 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.085 0.125 ;
END VIA45_FBD30_YEN

VIA VIA45_FBD30_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.125 0.085 0.025 ;
	LAYER VIA4 ;
		RECT 0.005 -0.115 0.055 0.015 ;
	LAYER M5 ;
		RECT -0.025 -0.125 0.085 0.025 ;
END VIA45_FBD30_YES

VIA VIA45_FBD30_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.085 -0.025 0.025 0.125 ;
	LAYER VIA4 ;
		RECT -0.055 -0.015 -0.005 0.115 ;
	LAYER M5 ;
		RECT -0.085 -0.025 0.025 0.125 ;
END VIA45_FBD30_YWN

VIA VIA45_FBD30_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.085 -0.125 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.055 -0.115 -0.005 0.015 ;
	LAYER M5 ;
		RECT -0.085 -0.125 0.025 0.025 ;
END VIA45_FBD30_YWS

VIA VIA45_PBDB_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.005 -0.045 0.165 0.045 ;
	LAYER VIA4 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA45_PBDB_E

VIA VIA45_PBDB_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.045 -0.005 0.045 0.165 ;
	LAYER VIA4 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA45_PBDB_N

VIA VIA45_PBDB_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.045 -0.165 0.045 0.005 ;
	LAYER VIA4 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M5 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA45_PBDB_S

VIA VIA45_PBDB_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.165 -0.045 0.005 0.045 ;
	LAYER VIA4 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M5 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA45_PBDB_W

VIA VIA45_PBDU_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.045 -0.025 0.165 0.025 ;
	LAYER VIA4 ;
		RECT -0.005 -0.025 0.125 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.045 0.145 0.045 ;
END VIA45_PBDU_E

VIA VIA45_PBDU_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.045 0.025 0.165 ;
	LAYER VIA4 ;
		RECT -0.025 -0.005 0.025 0.125 ;
	LAYER M5 ;
		RECT -0.045 -0.025 0.045 0.145 ;
END VIA45_PBDU_N

VIA VIA45_PBDU_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.165 0.025 0.045 ;
	LAYER VIA4 ;
		RECT -0.025 -0.125 0.025 0.005 ;
	LAYER M5 ;
		RECT -0.045 -0.145 0.045 0.025 ;
END VIA45_PBDU_S

VIA VIA45_PBDU_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.165 -0.025 0.045 0.025 ;
	LAYER VIA4 ;
		RECT -0.125 -0.025 0.005 0.025 ;
	LAYER M5 ;
		RECT -0.145 -0.045 0.025 0.045 ;
END VIA45_PBDU_W

VIA VIA45_PBDE_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.185 0.025 ;
	LAYER VIA4 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA45_PBDE_E

VIA VIA45_PBDE_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.025 0.185 ;
	LAYER VIA4 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA45_PBDE_N

VIA VIA45_PBDE_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.185 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M5 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA45_PBDE_S

VIA VIA45_PBDE_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M4 ;
		RECT -0.185 -0.025 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M5 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA45_PBDE_W

VIA VIA45_FBS25 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.05 -0.05 0.05 0.05 ;
END VIA45_FBS25

VIA VIA45_FBS25_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.025 0.075 0.075 ;
	LAYER VIA4 ;
		RECT 0 0 0.05 0.05 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.075 0.075 ;
END VIA45_FBS25_EN

VIA VIA45_FBS25_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.075 0.075 0.025 ;
	LAYER VIA4 ;
		RECT 0 -0.05 0.05 0 ;
	LAYER M5 ;
		RECT -0.025 -0.075 0.075 0.025 ;
END VIA45_FBS25_ES

VIA VIA45_FBS25_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.075 -0.025 0.025 0.075 ;
	LAYER VIA4 ;
		RECT -0.05 0 0 0.05 ;
	LAYER M5 ;
		RECT -0.075 -0.025 0.025 0.075 ;
END VIA45_FBS25_WN

VIA VIA45_FBS25_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.075 -0.075 0.025 0.025 ;
	LAYER VIA4 ;
		RECT -0.05 -0.05 0 0 ;
	LAYER M5 ;
		RECT -0.075 -0.075 0.025 0.025 ;
END VIA45_FBS25_WS

VIA VIA45_PBSU_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA45_PBSU_H

VIA VIA45_PBSU_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA45_PBSU_V

VIA VIA45_PBSB_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA45_PBSB_H

VIA VIA45_PBSB_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M4 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA4 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M5 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA45_PBSB_V


VIA VIA56_1cut DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA56_1cut

VIA VIA56_1cut_FAT_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.075 0.025 0.075 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.075 -0.025 0.075 0.025 ;
END VIA56_1cut_FAT_C

VIA VIA56_1cut_EN1415 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA56_1cut_EN1415

VIA VIA56_1stack_C DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.17 0.025 0.17 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA56_1stack_C

VIA VIA56_1stack_N DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.285 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA56_1stack_N

VIA VIA56_1stack_S DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.285 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA56_1stack_S

VIA VIA56_2cut_P1_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.155 ;
	LAYER VIA5 ;
		RECT -0.025 -0.015 0.025 0.115 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.125 ;
END VIA56_2cut_P1_N

VIA VIA56_2cut_P1_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.155 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.025 -0.115 0.025 0.015 ;
	LAYER M6 ;
		RECT -0.055 -0.125 0.055 0.025 ;
END VIA56_2cut_P1_S

VIA VIA56_2cut_P2_BLC DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.075 -0.055 0.075 0.055 ;
	LAYER VIA5 ;
		RECT -0.065 -0.025 0.065 0.025 ;
	LAYER M6 ;
		RECT -0.22 -0.025 0.22 0.025 ;
END VIA56_2cut_P2_BLC

VIA VIA56_2cut_P2_BLE DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA5 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M6 ;
		RECT -0.17 -0.025 0.27 0.025 ;
END VIA56_2cut_P2_BLE

VIA VIA56_2cut_P2_BLW DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M6 ;
		RECT -0.27 -0.025 0.17 0.025 ;
END VIA56_2cut_P2_BLW

VIA VIA56_2cut_P2_SLE DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA5 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M6 ;
		RECT -0.065 -0.025 0.375 0.025 ;
END VIA56_2cut_P2_SLE

VIA VIA56_2cut_P2_SLW DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M6 ;
		RECT -0.375 -0.025 0.065 0.025 ;
END VIA56_2cut_P2_SLW

VIA VIA56_2cut_P3_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.125 0.055 ;
	LAYER VIA5 ;
		RECT -0.015 -0.025 0.115 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.155 0.025 ;
END VIA56_2cut_P3_E

VIA VIA56_2cut_P3_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.125 -0.055 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.115 -0.025 0.015 0.025 ;
	LAYER M6 ;
		RECT -0.155 -0.025 0.055 0.025 ;
END VIA56_2cut_P3_W

VIA VIA56_4cut DEFAULT
	RESISTANCE 2.0000000000 ;
	LAYER M5 ;
		RECT -0.09 -0.12 0.09 0.12 ;
	LAYER VIA5 ;
		RECT -0.09 -0.09 -0.04 -0.04 ;
		RECT 0.04 -0.09 0.09 -0.04 ;
		RECT -0.09 0.04 -0.04 0.09 ;
		RECT 0.04 0.04 0.09 0.09 ;
	LAYER M6 ;
		RECT -0.12 -0.09 0.12 0.09 ;
END VIA56_4cut

VIA VIA56_FBD_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.165 0.085 ;
	LAYER VIA5 ;
		RECT 0.005 0.005 0.135 0.055 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.165 0.085 ;
END VIA56_FBD_XEN

VIA VIA56_FBD_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.085 0.165 0.025 ;
	LAYER VIA5 ;
		RECT 0.005 -0.055 0.135 -0.005 ;
	LAYER M6 ;
		RECT -0.025 -0.085 0.165 0.025 ;
END VIA56_FBD_XES

VIA VIA56_FBD_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.165 -0.025 0.025 0.085 ;
	LAYER VIA5 ;
		RECT -0.135 0.005 -0.005 0.055 ;
	LAYER M6 ;
		RECT -0.165 -0.025 0.025 0.085 ;
END VIA56_FBD_XWN

VIA VIA56_FBD_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.165 -0.085 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.135 -0.055 -0.005 -0.005 ;
	LAYER M6 ;
		RECT -0.165 -0.085 0.025 0.025 ;
END VIA56_FBD_XWS

VIA VIA56_FBD_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.085 0.165 ;
	LAYER VIA5 ;
		RECT 0.005 0.005 0.055 0.135 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.085 0.165 ;
END VIA56_FBD_YEN

VIA VIA56_FBD_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.165 0.085 0.025 ;
	LAYER VIA5 ;
		RECT 0.005 -0.135 0.055 -0.005 ;
	LAYER M6 ;
		RECT -0.025 -0.165 0.085 0.025 ;
END VIA56_FBD_YES

VIA VIA56_FBD_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.025 0.025 0.165 ;
	LAYER VIA5 ;
		RECT -0.055 0.005 -0.005 0.135 ;
	LAYER M6 ;
		RECT -0.085 -0.025 0.025 0.165 ;
END VIA56_FBD_YWN

VIA VIA56_FBD_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.165 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.055 -0.135 -0.005 -0.005 ;
	LAYER M6 ;
		RECT -0.085 -0.165 0.025 0.025 ;
END VIA56_FBD_YWS

VIA VIA56_FBS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.055 -0.055 0.055 0.055 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA56_FBS

VIA VIA56_FBS_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.085 0.085 ;
	LAYER VIA5 ;
		RECT 0.005 0.005 0.055 0.055 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.085 0.085 ;
END VIA56_FBS_EN

VIA VIA56_FBS_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.085 0.085 0.025 ;
	LAYER VIA5 ;
		RECT 0.005 -0.055 0.055 -0.005 ;
	LAYER M6 ;
		RECT -0.025 -0.085 0.085 0.025 ;
END VIA56_FBS_ES

VIA VIA56_FBS_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.025 0.025 0.085 ;
	LAYER VIA5 ;
		RECT -0.055 0.005 -0.005 0.055 ;
	LAYER M6 ;
		RECT -0.085 -0.025 0.025 0.085 ;
END VIA56_FBS_WN

VIA VIA56_FBS_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.085 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.055 -0.055 -0.005 -0.005 ;
	LAYER M6 ;
		RECT -0.085 -0.085 0.025 0.025 ;
END VIA56_FBS_WS

VIA VIA56_PBD_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.035 -0.025 0.175 0.025 ;
	LAYER VIA5 ;
		RECT 0.005 -0.025 0.135 0.025 ;
	LAYER M6 ;
		RECT -0.025 -0.055 0.165 0.055 ;
END VIA56_PBD_E

VIA VIA56_PBD_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.035 0.025 0.175 ;
	LAYER VIA5 ;
		RECT -0.025 0.005 0.025 0.135 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.165 ;
END VIA56_PBD_N

VIA VIA56_PBD_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.175 0.025 0.035 ;
	LAYER VIA5 ;
		RECT -0.025 -0.135 0.025 -0.005 ;
	LAYER M6 ;
		RECT -0.055 -0.165 0.055 0.025 ;
END VIA56_PBD_S

VIA VIA56_PBD_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.175 -0.025 0.035 0.025 ;
	LAYER VIA5 ;
		RECT -0.135 -0.025 -0.005 0.025 ;
	LAYER M6 ;
		RECT -0.165 -0.055 0.025 0.055 ;
END VIA56_PBD_W

VIA VIA56_PBS_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA56_PBS_H

VIA VIA56_PBS_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.055 0.055 0.055 ;
END VIA56_PBS_V

VIA VIA56_FBD20_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.145 0.065 ;
	LAYER VIA5 ;
		RECT -0.005 -0.005 0.125 0.045 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.145 0.065 ;
END VIA56_FBD20_XEN

VIA VIA56_FBD20_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.065 0.145 0.025 ;
	LAYER VIA5 ;
		RECT -0.005 -0.045 0.125 0.005 ;
	LAYER M6 ;
		RECT -0.025 -0.065 0.145 0.025 ;
END VIA56_FBD20_XES

VIA VIA56_FBD20_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.145 -0.025 0.025 0.065 ;
	LAYER VIA5 ;
		RECT -0.125 -0.005 0.005 0.045 ;
	LAYER M6 ;
		RECT -0.145 -0.025 0.025 0.065 ;
END VIA56_FBD20_XWN

VIA VIA56_FBD20_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.145 -0.065 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.125 -0.045 0.005 0.005 ;
	LAYER M6 ;
		RECT -0.145 -0.065 0.025 0.025 ;
END VIA56_FBD20_XWS

VIA VIA56_FBD20_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.065 0.145 ;
	LAYER VIA5 ;
		RECT -0.005 -0.005 0.045 0.125 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.065 0.145 ;
END VIA56_FBD20_YEN

VIA VIA56_FBD20_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.145 0.065 0.025 ;
	LAYER VIA5 ;
		RECT -0.005 -0.125 0.045 0.005 ;
	LAYER M6 ;
		RECT -0.025 -0.145 0.065 0.025 ;
END VIA56_FBD20_YES

VIA VIA56_FBD20_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.065 -0.025 0.025 0.145 ;
	LAYER VIA5 ;
		RECT -0.045 -0.005 0.005 0.125 ;
	LAYER M6 ;
		RECT -0.065 -0.025 0.025 0.145 ;
END VIA56_FBD20_YWN

VIA VIA56_FBD20_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.065 -0.145 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.045 -0.125 0.005 0.005 ;
	LAYER M6 ;
		RECT -0.065 -0.145 0.025 0.025 ;
END VIA56_FBD20_YWS

VIA VIA56_FBD30_XEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.125 0.085 ;
	LAYER VIA5 ;
		RECT -0.015 0.005 0.115 0.055 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.125 0.085 ;
END VIA56_FBD30_XEN

VIA VIA56_FBD30_XES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.085 0.125 0.025 ;
	LAYER VIA5 ;
		RECT -0.015 -0.055 0.115 -0.005 ;
	LAYER M6 ;
		RECT -0.025 -0.085 0.125 0.025 ;
END VIA56_FBD30_XES

VIA VIA56_FBD30_XWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.125 -0.025 0.025 0.085 ;
	LAYER VIA5 ;
		RECT -0.115 0.005 0.015 0.055 ;
	LAYER M6 ;
		RECT -0.125 -0.025 0.025 0.085 ;
END VIA56_FBD30_XWN

VIA VIA56_FBD30_XWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.125 -0.085 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.115 -0.055 0.015 -0.005 ;
	LAYER M6 ;
		RECT -0.125 -0.085 0.025 0.025 ;
END VIA56_FBD30_XWS

VIA VIA56_FBD30_YEN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.085 0.125 ;
	LAYER VIA5 ;
		RECT 0.005 -0.015 0.055 0.115 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.085 0.125 ;
END VIA56_FBD30_YEN

VIA VIA56_FBD30_YES DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.125 0.085 0.025 ;
	LAYER VIA5 ;
		RECT 0.005 -0.115 0.055 0.015 ;
	LAYER M6 ;
		RECT -0.025 -0.125 0.085 0.025 ;
END VIA56_FBD30_YES

VIA VIA56_FBD30_YWN DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.025 0.025 0.125 ;
	LAYER VIA5 ;
		RECT -0.055 -0.015 -0.005 0.115 ;
	LAYER M6 ;
		RECT -0.085 -0.025 0.025 0.125 ;
END VIA56_FBD30_YWN

VIA VIA56_FBD30_YWS DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.085 -0.125 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.055 -0.115 -0.005 0.015 ;
	LAYER M6 ;
		RECT -0.085 -0.125 0.025 0.025 ;
END VIA56_FBD30_YWS

VIA VIA56_PBDB_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.005 -0.045 0.165 0.045 ;
	LAYER VIA5 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA56_PBDB_E

VIA VIA56_PBDB_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.045 -0.005 0.045 0.165 ;
	LAYER VIA5 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA56_PBDB_N

VIA VIA56_PBDB_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.045 -0.165 0.045 0.005 ;
	LAYER VIA5 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M6 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA56_PBDB_S

VIA VIA56_PBDB_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.165 -0.045 0.005 0.045 ;
	LAYER VIA5 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M6 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA56_PBDB_W

VIA VIA56_PBDU_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.045 -0.025 0.165 0.025 ;
	LAYER VIA5 ;
		RECT -0.005 -0.025 0.125 0.025 ;
	LAYER M6 ;
		RECT -0.025 -0.045 0.145 0.045 ;
END VIA56_PBDU_E

VIA VIA56_PBDU_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.045 0.025 0.165 ;
	LAYER VIA5 ;
		RECT -0.025 -0.005 0.025 0.125 ;
	LAYER M6 ;
		RECT -0.045 -0.025 0.045 0.145 ;
END VIA56_PBDU_N

VIA VIA56_PBDU_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.165 0.025 0.045 ;
	LAYER VIA5 ;
		RECT -0.025 -0.125 0.025 0.005 ;
	LAYER M6 ;
		RECT -0.045 -0.145 0.045 0.025 ;
END VIA56_PBDU_S

VIA VIA56_PBDU_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.165 -0.025 0.045 0.025 ;
	LAYER VIA5 ;
		RECT -0.125 -0.025 0.005 0.025 ;
	LAYER M6 ;
		RECT -0.145 -0.045 0.025 0.045 ;
END VIA56_PBDU_W

VIA VIA56_PBDE_E DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.185 0.025 ;
	LAYER VIA5 ;
		RECT 0.015 -0.025 0.145 0.025 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.185 0.025 ;
END VIA56_PBDE_E

VIA VIA56_PBDE_N DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.025 0.185 ;
	LAYER VIA5 ;
		RECT -0.025 0.015 0.025 0.145 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.025 0.185 ;
END VIA56_PBDE_N

VIA VIA56_PBDE_S DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.185 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.025 -0.145 0.025 -0.015 ;
	LAYER M6 ;
		RECT -0.025 -0.185 0.025 0.025 ;
END VIA56_PBDE_S

VIA VIA56_PBDE_W DEFAULT
	RESISTANCE 4.5000000000 ;
	LAYER M5 ;
		RECT -0.185 -0.025 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.145 -0.025 -0.015 0.025 ;
	LAYER M6 ;
		RECT -0.185 -0.025 0.025 0.025 ;
END VIA56_PBDE_W

VIA VIA56_FBS25 DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
END VIA56_FBS25

VIA VIA56_FBS25_EN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.025 0.075 0.075 ;
	LAYER VIA5 ;
		RECT 0 0 0.05 0.05 ;
	LAYER M6 ;
		RECT -0.025 -0.025 0.075 0.075 ;
END VIA56_FBS25_EN

VIA VIA56_FBS25_ES DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.075 0.075 0.025 ;
	LAYER VIA5 ;
		RECT 0 -0.05 0.05 0 ;
	LAYER M6 ;
		RECT -0.025 -0.075 0.075 0.025 ;
END VIA56_FBS25_ES

VIA VIA56_FBS25_WN DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.075 -0.025 0.025 0.075 ;
	LAYER VIA5 ;
		RECT -0.05 0 0 0.05 ;
	LAYER M6 ;
		RECT -0.075 -0.025 0.025 0.075 ;
END VIA56_FBS25_WN

VIA VIA56_FBS25_WS DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.075 -0.075 0.025 0.025 ;
	LAYER VIA5 ;
		RECT -0.05 -0.05 0 0 ;
	LAYER M6 ;
		RECT -0.075 -0.075 0.025 0.025 ;
END VIA56_FBS25_WS

VIA VIA56_PBSU_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.055 -0.025 0.055 0.025 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.035 -0.05 0.035 0.05 ;
END VIA56_PBSU_H

VIA VIA56_PBSU_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.025 -0.055 0.025 0.055 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.05 -0.035 0.05 0.035 ;
END VIA56_PBSU_V

VIA VIA56_PBSB_H DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.05 -0.035 0.05 0.035 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.025 -0.055 0.025 0.055 ;
END VIA56_PBSB_H

VIA VIA56_PBSB_V DEFAULT
	RESISTANCE 8.0000000000 ;
	LAYER M5 ;
		RECT -0.035 -0.05 0.035 0.05 ;
	LAYER VIA5 ;
		RECT -0.025 -0.025 0.025 0.025 ;
	LAYER M6 ;
		RECT -0.055 -0.025 0.055 0.025 ;
END VIA56_PBSB_V


VIA VIA67_1cut DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.09 -0.065 0.09 0.065 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.09 ;
END VIA67_1cut

VIA VIA67_1cut_FAT_C DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.115 -0.065 0.115 0.065 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.05 -0.115 0.05 0.115 ;
END VIA67_1cut_FAT_C

VIA VIA67_1cut_FAT_H DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.115 -0.065 0.115 0.065 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.115 -0.05 0.115 0.05 ;
END VIA67_1cut_FAT_H

VIA VIA67_1cut_FAT_V DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.065 -0.115 0.065 0.115 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.05 -0.115 0.05 0.115 ;
END VIA67_1cut_FAT_V

VIA VIA67_1cut_H DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.09 -0.065 0.09 0.065 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.09 -0.05 0.09 0.05 ;
END VIA67_1cut_H

VIA VIA67_1cut_V DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.065 -0.09 0.065 0.09 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.09 ;
END VIA67_1cut_V

VIA VIA67_2cut_P1_E DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.09 -0.065 0.29 0.065 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT 0.15 -0.05 0.25 0.05 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.25 0.09 ;
END VIA67_2cut_P1_E

VIA VIA67_2cut_P1_N DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.065 -0.09 0.065 0.29 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT -0.05 0.15 0.05 0.25 ;
	LAYER M7 ;
		RECT -0.09 -0.05 0.09 0.25 ;
END VIA67_2cut_P1_N

VIA VIA67_2cut_P1_S DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.065 -0.29 0.065 0.09 ;
	LAYER VIA6 ;
		RECT -0.05 -0.25 0.05 -0.15 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.09 -0.25 0.09 0.05 ;
END VIA67_2cut_P1_S

VIA VIA67_2cut_P1_W DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.29 -0.065 0.09 0.065 ;
	LAYER VIA6 ;
		RECT -0.25 -0.05 -0.15 0.05 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.25 -0.09 0.05 0.09 ;
END VIA67_2cut_P1_W

VIA VIA67_2cut_P3_E DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.065 -0.09 0.265 0.09 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT 0.15 -0.05 0.25 0.05 ;
	LAYER M7 ;
		RECT -0.09 -0.05 0.29 0.05 ;
END VIA67_2cut_P3_E

VIA VIA67_2cut_P3_N DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.09 -0.065 0.09 0.265 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT -0.05 0.15 0.05 0.25 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.29 ;
END VIA67_2cut_P3_N

VIA VIA67_2cut_P3_S DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.09 -0.265 0.09 0.065 ;
	LAYER VIA6 ;
		RECT -0.05 -0.25 0.05 -0.15 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.05 -0.29 0.05 0.09 ;
END VIA67_2cut_P3_S

VIA VIA67_2cut_P3_W DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.265 -0.09 0.065 0.09 ;
	LAYER VIA6 ;
		RECT -0.25 -0.05 -0.15 0.05 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.29 -0.05 0.09 0.05 ;
END VIA67_2cut_P3_W

VIA VIA67_4cut DEFAULT
	RESISTANCE 0.6250000000 ;
	LAYER M6 ;
		RECT -0.205 -0.18 0.205 0.18 ;
	LAYER VIA6 ;
		RECT -0.165 -0.165 -0.065 -0.065 ;
		RECT 0.065 -0.165 0.165 -0.065 ;
		RECT -0.165 0.065 -0.065 0.165 ;
		RECT 0.065 0.065 0.165 0.165 ;
	LAYER M7 ;
		RECT -0.165 -0.205 0.165 0.205 ;
END VIA67_4cut

VIA VIA67_FBD_XEN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.05 -0.05 0.33 0.13 ;
	LAYER VIA6 ;
		RECT -0.01 -0.01 0.09 0.09 ;
		RECT 0.19 -0.01 0.29 0.09 ;
	LAYER M7 ;
		RECT -0.05 -0.05 0.33 0.13 ;
END VIA67_FBD_XEN

VIA VIA67_FBD_XES DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.05 -0.13 0.33 0.05 ;
	LAYER VIA6 ;
		RECT -0.01 -0.09 0.09 0.01 ;
		RECT 0.19 -0.09 0.29 0.01 ;
	LAYER M7 ;
		RECT -0.05 -0.13 0.33 0.05 ;
END VIA67_FBD_XES

VIA VIA67_FBD_XWN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.33 -0.05 0.05 0.13 ;
	LAYER VIA6 ;
		RECT -0.29 -0.01 -0.19 0.09 ;
		RECT -0.09 -0.01 0.01 0.09 ;
	LAYER M7 ;
		RECT -0.33 -0.05 0.05 0.13 ;
END VIA67_FBD_XWN

VIA VIA67_FBD_XWS DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.33 -0.13 0.05 0.05 ;
	LAYER VIA6 ;
		RECT -0.29 -0.09 -0.19 0.01 ;
		RECT -0.09 -0.09 0.01 0.01 ;
	LAYER M7 ;
		RECT -0.33 -0.13 0.05 0.05 ;
END VIA67_FBD_XWS

VIA VIA67_FBD_YEN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.05 -0.05 0.13 0.33 ;
	LAYER VIA6 ;
		RECT -0.01 -0.01 0.09 0.09 ;
		RECT -0.01 0.19 0.09 0.29 ;
	LAYER M7 ;
		RECT -0.05 -0.05 0.13 0.33 ;
END VIA67_FBD_YEN

VIA VIA67_FBD_YES DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.05 -0.33 0.13 0.05 ;
	LAYER VIA6 ;
		RECT -0.01 -0.29 0.09 -0.19 ;
		RECT -0.01 -0.09 0.09 0.01 ;
	LAYER M7 ;
		RECT -0.05 -0.33 0.13 0.05 ;
END VIA67_FBD_YES

VIA VIA67_FBD_YWN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.13 -0.05 0.05 0.33 ;
	LAYER VIA6 ;
		RECT -0.09 -0.01 0.01 0.09 ;
		RECT -0.09 0.19 0.01 0.29 ;
	LAYER M7 ;
		RECT -0.13 -0.05 0.05 0.33 ;
END VIA67_FBD_YWN

VIA VIA67_FBD_YWS DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M6 ;
		RECT -0.13 -0.33 0.05 0.05 ;
	LAYER VIA6 ;
		RECT -0.09 -0.29 0.01 -0.19 ;
		RECT -0.09 -0.09 0.01 0.01 ;
	LAYER M7 ;
		RECT -0.13 -0.33 0.05 0.05 ;
END VIA67_FBD_YWS

VIA VIA67_FBS DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.09 -0.09 0.09 0.09 ;
	LAYER VIA6 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M7 ;
		RECT -0.09 -0.09 0.09 0.09 ;
END VIA67_FBS

VIA VIA67_FBS_EN DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.05 -0.05 0.13 0.13 ;
	LAYER VIA6 ;
		RECT -0.01 -0.01 0.09 0.09 ;
	LAYER M7 ;
		RECT -0.05 -0.05 0.13 0.13 ;
END VIA67_FBS_EN

VIA VIA67_FBS_ES DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.05 -0.13 0.13 0.05 ;
	LAYER VIA6 ;
		RECT -0.01 -0.09 0.09 0.01 ;
	LAYER M7 ;
		RECT -0.05 -0.13 0.13 0.05 ;
END VIA67_FBS_ES

VIA VIA67_FBS_WN DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.13 -0.05 0.05 0.13 ;
	LAYER VIA6 ;
		RECT -0.09 -0.01 0.01 0.09 ;
	LAYER M7 ;
		RECT -0.13 -0.05 0.05 0.13 ;
END VIA67_FBS_WN

VIA VIA67_FBS_WS DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M6 ;
		RECT -0.13 -0.13 0.05 0.05 ;
	LAYER VIA6 ;
		RECT -0.09 -0.09 0.01 0.01 ;
	LAYER M7 ;
		RECT -0.13 -0.13 0.05 0.05 ;
END VIA67_FBS_WS


VIA VIA78_1cut DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.09 0.05 ;
END VIA78_1cut

VIA VIA78_1cut_FAT_C DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.115 0.05 0.115 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.115 -0.05 0.115 0.05 ;
END VIA78_1cut_FAT_C

VIA VIA78_1cut_FAT_H DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.115 -0.05 0.115 0.05 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.115 -0.05 0.115 0.05 ;
END VIA78_1cut_FAT_H

VIA VIA78_1cut_FAT_V DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.115 0.05 0.115 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.05 -0.115 0.05 0.115 ;
END VIA78_1cut_FAT_V

VIA VIA78_1cut_H DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.09 -0.05 0.09 0.05 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.09 0.05 ;
END VIA78_1cut_H

VIA VIA78_1cut_V DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.05 -0.09 0.05 0.09 ;
END VIA78_1cut_V

VIA VIA78_1stack_N DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.43 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.09 0.05 ;
END VIA78_1stack_N

VIA VIA78_1stack_S DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.43 0.05 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.09 0.05 ;
END VIA78_1stack_S

VIA VIA78_2cut_P1_E DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.09 -0.05 0.29 0.05 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT 0.15 -0.05 0.25 0.05 ;
	LAYER M8 ;
		RECT -0.05 -0.09 0.25 0.09 ;
END VIA78_2cut_P1_E

VIA VIA78_2cut_P1_N DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.29 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT -0.05 0.15 0.05 0.25 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.09 0.25 ;
END VIA78_2cut_P1_N

VIA VIA78_2cut_P1_S DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.29 0.05 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.25 0.05 -0.15 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.25 0.09 0.05 ;
END VIA78_2cut_P1_S

VIA VIA78_2cut_P1_W DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.29 -0.05 0.09 0.05 ;
	LAYER VIA7 ;
		RECT -0.25 -0.05 -0.15 0.05 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.25 -0.09 0.05 0.09 ;
END VIA78_2cut_P1_W

VIA VIA78_2cut_P3_E DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.25 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT 0.15 -0.05 0.25 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.29 0.05 ;
END VIA78_2cut_P3_E

VIA VIA78_2cut_P3_N DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.09 -0.05 0.09 0.25 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT -0.05 0.15 0.05 0.25 ;
	LAYER M8 ;
		RECT -0.05 -0.09 0.05 0.29 ;
END VIA78_2cut_P3_N

VIA VIA78_2cut_P3_S DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.09 -0.25 0.09 0.05 ;
	LAYER VIA7 ;
		RECT -0.05 -0.25 0.05 -0.15 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.05 -0.29 0.05 0.09 ;
END VIA78_2cut_P3_S

VIA VIA78_2cut_P3_W DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.25 -0.09 0.05 0.09 ;
	LAYER VIA7 ;
		RECT -0.25 -0.05 -0.15 0.05 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.29 -0.05 0.09 0.05 ;
END VIA78_2cut_P3_W

VIA VIA78_4cut DEFAULT
	RESISTANCE 0.6250000000 ;
	LAYER M7 ;
		RECT -0.165 -0.205 0.165 0.205 ;
	LAYER VIA7 ;
		RECT -0.165 -0.165 -0.065 -0.065 ;
		RECT 0.065 -0.165 0.165 -0.065 ;
		RECT -0.165 0.065 -0.065 0.165 ;
		RECT 0.065 0.065 0.165 0.165 ;
	LAYER M8 ;
		RECT -0.205 -0.165 0.205 0.165 ;
END VIA78_4cut

VIA VIA78_2stack_N DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.09 0.05 0.43 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
		RECT -0.05 0.15 0.05 0.25 ;
	LAYER M8 ;
		RECT -0.09 -0.05 0.09 0.25 ;
END VIA78_2stack_N

VIA VIA78_2stack_S DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.43 0.05 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.25 0.05 -0.15 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.25 0.09 0.05 ;
END VIA78_2stack_S

VIA VIA78_FBD_XEN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.05 0.33 0.13 ;
	LAYER VIA7 ;
		RECT -0.01 -0.01 0.09 0.09 ;
		RECT 0.19 -0.01 0.29 0.09 ;
	LAYER M8 ;
		RECT -0.05 -0.05 0.33 0.13 ;
END VIA78_FBD_XEN

VIA VIA78_FBD_XES DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.13 0.33 0.05 ;
	LAYER VIA7 ;
		RECT -0.01 -0.09 0.09 0.01 ;
		RECT 0.19 -0.09 0.29 0.01 ;
	LAYER M8 ;
		RECT -0.05 -0.13 0.33 0.05 ;
END VIA78_FBD_XES

VIA VIA78_FBD_XWN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.33 -0.05 0.05 0.13 ;
	LAYER VIA7 ;
		RECT -0.29 -0.01 -0.19 0.09 ;
		RECT -0.09 -0.01 0.01 0.09 ;
	LAYER M8 ;
		RECT -0.33 -0.05 0.05 0.13 ;
END VIA78_FBD_XWN

VIA VIA78_FBD_XWS DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.33 -0.13 0.05 0.05 ;
	LAYER VIA7 ;
		RECT -0.29 -0.09 -0.19 0.01 ;
		RECT -0.09 -0.09 0.01 0.01 ;
	LAYER M8 ;
		RECT -0.33 -0.13 0.05 0.05 ;
END VIA78_FBD_XWS

VIA VIA78_FBD_YEN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.05 0.13 0.33 ;
	LAYER VIA7 ;
		RECT -0.01 -0.01 0.09 0.09 ;
		RECT -0.01 0.19 0.09 0.29 ;
	LAYER M8 ;
		RECT -0.05 -0.05 0.13 0.33 ;
END VIA78_FBD_YEN

VIA VIA78_FBD_YES DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.05 -0.33 0.13 0.05 ;
	LAYER VIA7 ;
		RECT -0.01 -0.29 0.09 -0.19 ;
		RECT -0.01 -0.09 0.09 0.01 ;
	LAYER M8 ;
		RECT -0.05 -0.33 0.13 0.05 ;
END VIA78_FBD_YES

VIA VIA78_FBD_YWN DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.13 -0.05 0.05 0.33 ;
	LAYER VIA7 ;
		RECT -0.09 -0.01 0.01 0.09 ;
		RECT -0.09 0.19 0.01 0.29 ;
	LAYER M8 ;
		RECT -0.13 -0.05 0.05 0.33 ;
END VIA78_FBD_YWN

VIA VIA78_FBD_YWS DEFAULT
	RESISTANCE 1.2500000000 ;
	LAYER M7 ;
		RECT -0.13 -0.33 0.05 0.05 ;
	LAYER VIA7 ;
		RECT -0.09 -0.29 0.01 -0.19 ;
		RECT -0.09 -0.09 0.01 0.01 ;
	LAYER M8 ;
		RECT -0.13 -0.33 0.05 0.05 ;
END VIA78_FBD_YWS

VIA VIA78_FBS DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.09 -0.09 0.09 0.09 ;
	LAYER VIA7 ;
		RECT -0.05 -0.05 0.05 0.05 ;
	LAYER M8 ;
		RECT -0.09 -0.09 0.09 0.09 ;
END VIA78_FBS

VIA VIA78_FBS_EN DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.05 0.13 0.13 ;
	LAYER VIA7 ;
		RECT -0.01 -0.01 0.09 0.09 ;
	LAYER M8 ;
		RECT -0.05 -0.05 0.13 0.13 ;
END VIA78_FBS_EN

VIA VIA78_FBS_ES DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.05 -0.13 0.13 0.05 ;
	LAYER VIA7 ;
		RECT -0.01 -0.09 0.09 0.01 ;
	LAYER M8 ;
		RECT -0.05 -0.13 0.13 0.05 ;
END VIA78_FBS_ES

VIA VIA78_FBS_WN DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.13 -0.05 0.05 0.13 ;
	LAYER VIA7 ;
		RECT -0.09 -0.01 0.01 0.09 ;
	LAYER M8 ;
		RECT -0.13 -0.05 0.05 0.13 ;
END VIA78_FBS_WN

VIA VIA78_FBS_WS DEFAULT
	RESISTANCE 2.5000000000 ;
	LAYER M7 ;
		RECT -0.13 -0.13 0.05 0.05 ;
	LAYER VIA7 ;
		RECT -0.09 -0.09 0.01 0.01 ;
	LAYER M8 ;
		RECT -0.13 -0.13 0.05 0.05 ;
END VIA78_FBS_WS


VIA VIA89_1cut DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M8 ;
		RECT -0.26 -0.2 0.26 0.2 ;
	LAYER VIA8 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 0.26 ;
END VIA89_1cut

VIA VIA89_1cut_H DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M8 ;
		RECT -0.26 -0.2 0.26 0.2 ;
	LAYER VIA8 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M9 ;
		RECT -0.26 -0.2 0.26 0.2 ;
END VIA89_1cut_H

VIA VIA89_1cut_V DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M8 ;
		RECT -0.2 -0.26 0.2 0.26 ;
	LAYER VIA8 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 0.26 ;
END VIA89_1cut_V

VIA VIA89_2cut_P1_E DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M8 ;
		RECT -0.26 -0.2 0.96 0.2 ;
	LAYER VIA8 ;
		RECT -0.18 -0.18 0.18 0.18 ;
		RECT 0.52 -0.18 0.88 0.18 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.9 0.26 ;
END VIA89_2cut_P1_E

VIA VIA89_2cut_P1_W DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M8 ;
		RECT -0.96 -0.2 0.26 0.2 ;
	LAYER VIA8 ;
		RECT -0.88 -0.18 -0.52 0.18 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M9 ;
		RECT -0.9 -0.26 0.2 0.26 ;
END VIA89_2cut_P1_W

VIA VIA89_2cut_P3_N DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M8 ;
		RECT -0.26 -0.2 0.26 0.9 ;
	LAYER VIA8 ;
		RECT -0.18 -0.18 0.18 0.18 ;
		RECT -0.18 0.52 0.18 0.88 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 0.96 ;
END VIA89_2cut_P3_N

VIA VIA89_2cut_P3_S DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M8 ;
		RECT -0.26 -0.9 0.26 0.2 ;
	LAYER VIA8 ;
		RECT -0.18 -0.88 0.18 -0.52 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M9 ;
		RECT -0.2 -0.96 0.2 0.26 ;
END VIA89_2cut_P3_S

VIA VIA89_4cut DEFAULT
	RESISTANCE 0.0675000000 ;
	LAYER M8 ;
		RECT -0.71 -0.65 0.71 0.65 ;
	LAYER VIA8 ;
		RECT -0.63 -0.63 -0.27 -0.27 ;
		RECT 0.27 -0.63 0.63 -0.27 ;
		RECT -0.63 0.27 -0.27 0.63 ;
		RECT 0.27 0.27 0.63 0.63 ;
	LAYER M9 ;
		RECT -0.65 -0.71 0.65 0.71 ;
END VIA89_4cut

VIA VIA89_FBS DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M8 ;
		RECT -0.26 -0.26 0.26 0.26 ;
	LAYER VIA8 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M9 ;
		RECT -0.26 -0.26 0.26 0.26 ;
END VIA89_FBS


VIA VIA910_1cut DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.26 0.2 ;
END VIA910_1cut

VIA VIA910_1cut_H DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M9 ;
		RECT -0.26 -0.2 0.26 0.2 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.26 0.2 ;
END VIA910_1cut_H

VIA VIA910_1cut_V DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.2 -0.26 0.2 0.26 ;
END VIA910_1cut_V

VIA VIA910_1stack_N DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 1.155 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.26 0.2 ;
END VIA910_1stack_N

VIA VIA910_1stack_S DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M9 ;
		RECT -0.2 -1.155 0.2 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.26 0.2 ;
END VIA910_1stack_S

VIA VIA910_2cut_P3_E DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.9 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
		RECT 0.52 -0.18 0.88 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.96 0.2 ;
END VIA910_2cut_P3_E

VIA VIA910_2cut_P3_W DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M9 ;
		RECT -0.9 -0.26 0.2 0.26 ;
	LAYER VIA9 ;
		RECT -0.88 -0.18 -0.52 0.18 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.96 -0.2 0.26 0.2 ;
END VIA910_2cut_P3_W

VIA VIA910_2cut_P1_N DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 0.96 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
		RECT -0.18 0.52 0.18 0.88 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.26 0.9 ;
END VIA910_2cut_P1_N

VIA VIA910_2cut_P1_S DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M9 ;
		RECT -0.2 -0.96 0.2 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.88 0.18 -0.52 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.9 0.26 0.2 ;
END VIA910_2cut_P1_S

VIA VIA910_2stack_N DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M9 ;
		RECT -0.2 -0.26 0.2 1.155 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
		RECT -0.18 0.52 0.18 0.88 ;
	LAYER M10 ;
		RECT -0.26 -0.2 0.26 0.9 ;
END VIA910_2stack_N

VIA VIA910_2stack_S DEFAULT
	RESISTANCE 0.1350000000 ;
	LAYER M9 ;
		RECT -0.2 -1.155 0.2 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.88 0.18 -0.52 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.9 0.26 0.2 ;
END VIA910_2stack_S

VIA VIA910_4cut DEFAULT
	RESISTANCE 0.0675000000 ;
	LAYER M9 ;
		RECT -0.65 -0.71 0.65 0.71 ;
	LAYER VIA9 ;
		RECT -0.63 -0.63 -0.27 -0.27 ;
		RECT 0.27 -0.63 0.63 -0.27 ;
		RECT -0.63 0.27 -0.27 0.63 ;
		RECT 0.27 0.27 0.63 0.63 ;
	LAYER M10 ;
		RECT -0.71 -0.65 0.71 0.65 ;
END VIA910_4cut

VIA VIA910_FBS DEFAULT
	RESISTANCE 0.2700000000 ;
	LAYER M9 ;
		RECT -0.26 -0.26 0.26 0.26 ;
	LAYER VIA9 ;
		RECT -0.18 -0.18 0.18 0.18 ;
	LAYER M10 ;
		RECT -0.26 -0.26 0.26 0.26 ;
END VIA910_FBS


VIA VIA10AP_1cut DEFAULT
	RESISTANCE 0.0640000000 ;
	LAYER M10 ;
		RECT -2 -2 2 2 ;
	LAYER RV ;
		RECT -1.5 -1.5 1.5 1.5 ;
	LAYER AP ;
		RECT -2 -2 2 2 ;
END VIA10AP_1cut

### RV 2um x 2um is only allowed in plymide process, if below device is turn on, please turn off above.
#VIA VIA10AP_1cut DEFAULT
#	RESISTANCE 0.0640000000 ;
#	LAYER M10 ;
#		RECT -1.5 -1.5 1.5 1.5 ;
#	LAYER RV ;
#		RECT -1 -1 1 1 ;
#	LAYER AP ;
#		RECT -1.5 -1.5 1.5 1.5 ;
#END VIA10AP_1cut


VIARULE VIAGEN12 GENERATE
    LAYER M1 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER M2 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER VIA1 ;
        RECT -0.025 -0.025 0.025 0.025 ;
        SPACING 0.13 BY 0.13 ;
END VIAGEN12


VIARULE VIAGEN12_RECT GENERATE
    LAYER M1 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER M2 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER VIA1 ;
        RECT -0.025000 -0.025000 0.105000 0.025000 ;
        SPACING 0.210000 BY 0.130000 ;
END VIAGEN12_RECT


VIARULE VIAGEN23 GENERATE
    LAYER M2 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER M3 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER VIA2 ;
        RECT -0.025 -0.025 0.025 0.025 ;
        SPACING 0.13 BY 0.13 ;
END VIAGEN23


VIARULE VIAGEN23_RECT GENERATE
    LAYER M2 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER M3 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER VIA2 ;
        RECT -0.025000 -0.025000 0.105000 0.025000 ;
        SPACING 0.210000 BY 0.130000 ;
END VIAGEN23_RECT


VIARULE VIAGEN34 GENERATE
    LAYER M3 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER M4 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER VIA3 ;
        RECT -0.025 -0.025 0.025 0.025 ;
        SPACING 0.13 BY 0.13 ;
END VIAGEN34


VIARULE VIAGEN34_RECT GENERATE
    LAYER M3 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER M4 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER VIA3 ;
        RECT -0.025000 -0.025000 0.105000 0.025000 ;
        SPACING 0.210000 BY 0.130000 ;
END VIAGEN34_RECT


VIARULE VIAGEN45 GENERATE
    LAYER M4 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER M5 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER VIA4 ;
        RECT -0.025 -0.025 0.025 0.025 ;
        SPACING 0.13 BY 0.13 ;
END VIAGEN45


VIARULE VIAGEN45_RECT GENERATE
    LAYER M4 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER M5 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER VIA4 ;
        RECT -0.025000 -0.025000 0.105000 0.025000 ;
        SPACING 0.210000 BY 0.130000 ;
END VIAGEN45_RECT


VIARULE VIAGEN56 GENERATE
    LAYER M5 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER M6 ;
        ENCLOSURE 0.03 0 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER VIA5 ;
        RECT -0.025 -0.025 0.025 0.025 ;
        SPACING 0.13 BY 0.13 ;
END VIAGEN56


VIARULE VIAGEN56_RECT GENERATE
    LAYER M5 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER M6 ;
        ENCLOSURE 0.040000 0.000000 ;
        WIDTH 0.050000 TO 4.500000 ;
    LAYER VIA5 ;
        RECT -0.025000 -0.025000 0.105000 0.025000 ;
        SPACING 0.210000 BY 0.130000 ;
END VIAGEN56_RECT


VIARULE VIAGEN67 GENERATE
    LAYER M6 ;
        ENCLOSURE 0.04 0.015 ;
        WIDTH 0.05 TO 4.5 ;
    LAYER M7 ;
        ENCLOSURE 0.04 0 ;
        WIDTH 0.1 TO 12 ;
    LAYER VIA6 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        SPACING 0.23 BY 0.23 ;
END VIAGEN67


VIARULE VIAGEN78 GENERATE
    LAYER M7 ;
        ENCLOSURE 0.04 0 ;
        WIDTH 0.1 TO 12 ;
    LAYER M8 ;
        ENCLOSURE 0.04 0 ;
        WIDTH 0.1 TO 12 ;
    LAYER VIA7 ;
        RECT -0.05 -0.05 0.05 0.05 ;
        SPACING 0.23 BY 0.23 ;
END VIAGEN78


VIARULE VIAGEN89 GENERATE
    LAYER M8 ;
        ENCLOSURE 0.08 0.02 ;
        WIDTH 0.1 TO 12 ;
    LAYER M9 ;
        ENCLOSURE 0.08 0.02 ;
        WIDTH 0.4 TO 12 ;
    LAYER VIA8 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.9 BY 0.9 ;
END VIAGEN89


VIARULE VIAGEN910 GENERATE
    LAYER M9 ;
        ENCLOSURE 0.08 0.02 ;
        WIDTH 0.4 TO 12 ;
    LAYER M10 ;
        ENCLOSURE 0.08 0.02 ;
        WIDTH 0.4 TO 12 ;
    LAYER VIA9 ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.9 BY 0.9 ;
END VIAGEN910


VIARULE VIAGEN10AP GENERATE
    LAYER M10 ;
        ENCLOSURE 0.500000 0.500000 ;
        WIDTH 0.4 TO 12 ;
    LAYER AP ;
        ENCLOSURE 0.500000 0.500000 ;
        WIDTH 2.000000 TO 35.000000 ;
    LAYER RV ;
        RECT -1.500000 -1.500000 1.500000 1.500000 ;
        SPACING 5.000000 BY 5.000000 ;
END VIAGEN10AP

### RV 2um x 2um is only allowed in plymide process, if below VIARULE is turn on, please turn off above
#VIARULE VIAGEN10AP GENERATE
#    LAYER M10 ;
#        ENCLOSURE 0.500000 0.500000 ;
#        WIDTH 0.4 TO 12 ;
#    LAYER AP ;
#        ENCLOSURE 0.500000 0.500000 ;
#        WIDTH 2.000000 TO 35.000000 ;
#    LAYER RV ;
#        RECT -1.000000 -1.000000 1.000000 1.000000 ;
#        SPACING 4.000000 BY 4.000000 ;
#END VIAGEN10AP

