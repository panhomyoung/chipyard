module mem_ext(
  input  [8:0]  RW0_addr,
  input         RW0_clk,
  input  [63:0] RW0_wdata,
  output [63:0] RW0_rdata,
  input         RW0_en,
  input         RW0_wmode,
  input  [7:0]  RW0_wmask
);
  wire [8:0] mem_0_0_0_RW0_addr;
  wire  mem_0_0_0_RW0_clk;
  wire [7:0] mem_0_0_0_RW0_wdata;
  wire [7:0] mem_0_0_0_RW0_rdata;
  wire  mem_0_0_0_RW0_en;
  wire  mem_0_0_0_RW0_wmode;
  wire  mem_0_0_0_RW0_wmask;
  wire [8:0] mem_0_1_0_RW0_addr;
  wire  mem_0_1_0_RW0_clk;
  wire [7:0] mem_0_1_0_RW0_wdata;
  wire [7:0] mem_0_1_0_RW0_rdata;
  wire  mem_0_1_0_RW0_en;
  wire  mem_0_1_0_RW0_wmode;
  wire  mem_0_1_0_RW0_wmask;
  wire [8:0] mem_0_2_0_RW0_addr;
  wire  mem_0_2_0_RW0_clk;
  wire [7:0] mem_0_2_0_RW0_wdata;
  wire [7:0] mem_0_2_0_RW0_rdata;
  wire  mem_0_2_0_RW0_en;
  wire  mem_0_2_0_RW0_wmode;
  wire  mem_0_2_0_RW0_wmask;
  wire [8:0] mem_0_3_0_RW0_addr;
  wire  mem_0_3_0_RW0_clk;
  wire [7:0] mem_0_3_0_RW0_wdata;
  wire [7:0] mem_0_3_0_RW0_rdata;
  wire  mem_0_3_0_RW0_en;
  wire  mem_0_3_0_RW0_wmode;
  wire  mem_0_3_0_RW0_wmask;
  wire [8:0] mem_0_4_0_RW0_addr;
  wire  mem_0_4_0_RW0_clk;
  wire [7:0] mem_0_4_0_RW0_wdata;
  wire [7:0] mem_0_4_0_RW0_rdata;
  wire  mem_0_4_0_RW0_en;
  wire  mem_0_4_0_RW0_wmode;
  wire  mem_0_4_0_RW0_wmask;
  wire [8:0] mem_0_5_0_RW0_addr;
  wire  mem_0_5_0_RW0_clk;
  wire [7:0] mem_0_5_0_RW0_wdata;
  wire [7:0] mem_0_5_0_RW0_rdata;
  wire  mem_0_5_0_RW0_en;
  wire  mem_0_5_0_RW0_wmode;
  wire  mem_0_5_0_RW0_wmask;
  wire [8:0] mem_0_6_0_RW0_addr;
  wire  mem_0_6_0_RW0_clk;
  wire [7:0] mem_0_6_0_RW0_wdata;
  wire [7:0] mem_0_6_0_RW0_rdata;
  wire  mem_0_6_0_RW0_en;
  wire  mem_0_6_0_RW0_wmode;
  wire  mem_0_6_0_RW0_wmask;
  wire [8:0] mem_0_7_0_RW0_addr;
  wire  mem_0_7_0_RW0_clk;
  wire [7:0] mem_0_7_0_RW0_wdata;
  wire [7:0] mem_0_7_0_RW0_rdata;
  wire  mem_0_7_0_RW0_en;
  wire  mem_0_7_0_RW0_wmode;
  wire  mem_0_7_0_RW0_wmask;
  wire [7:0] RW0_rdata_0_0_0 = mem_0_0_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_1_0 = mem_0_1_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_2_0 = mem_0_2_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_3_0 = mem_0_3_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_4_0 = mem_0_4_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_5_0 = mem_0_5_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_6_0 = mem_0_6_0_RW0_rdata;
  wire [7:0] RW0_rdata_0_7_0 = mem_0_7_0_RW0_rdata;
  wire [15:0] _GEN_0 = {RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [23:0] _GEN_1 = {RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [31:0] _GEN_2 = {RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [39:0] _GEN_3 = {RW0_rdata_0_4_0,RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [47:0] _GEN_4 = {RW0_rdata_0_5_0,RW0_rdata_0_4_0,RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0}
    ;
  wire [55:0] _GEN_5 = {RW0_rdata_0_6_0,RW0_rdata_0_5_0,RW0_rdata_0_4_0,RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,
    RW0_rdata_0_0_0};
  wire [63:0] RW0_rdata_0_0 = {RW0_rdata_0_7_0,RW0_rdata_0_6_0,RW0_rdata_0_5_0,RW0_rdata_0_4_0,RW0_rdata_0_3_0,
    RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [15:0] _GEN_6 = {RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [23:0] _GEN_7 = {RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [31:0] _GEN_8 = {RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [39:0] _GEN_9 = {RW0_rdata_0_4_0,RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0};
  wire [47:0] _GEN_10 = {RW0_rdata_0_5_0,RW0_rdata_0_4_0,RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0,RW0_rdata_0_0_0
    };
  wire [55:0] _GEN_11 = {RW0_rdata_0_6_0,RW0_rdata_0_5_0,RW0_rdata_0_4_0,RW0_rdata_0_3_0,RW0_rdata_0_2_0,RW0_rdata_0_1_0
    ,RW0_rdata_0_0_0};
  split_mem_ext mem_0_0_0 (
    .RW0_addr(mem_0_0_0_RW0_addr),
    .RW0_clk(mem_0_0_0_RW0_clk),
    .RW0_wdata(mem_0_0_0_RW0_wdata),
    .RW0_rdata(mem_0_0_0_RW0_rdata),
    .RW0_en(mem_0_0_0_RW0_en),
    .RW0_wmode(mem_0_0_0_RW0_wmode),
    .RW0_wmask(mem_0_0_0_RW0_wmask)
  );
  split_mem_ext mem_0_1_0 (
    .RW0_addr(mem_0_1_0_RW0_addr),
    .RW0_clk(mem_0_1_0_RW0_clk),
    .RW0_wdata(mem_0_1_0_RW0_wdata),
    .RW0_rdata(mem_0_1_0_RW0_rdata),
    .RW0_en(mem_0_1_0_RW0_en),
    .RW0_wmode(mem_0_1_0_RW0_wmode),
    .RW0_wmask(mem_0_1_0_RW0_wmask)
  );
  split_mem_ext mem_0_2_0 (
    .RW0_addr(mem_0_2_0_RW0_addr),
    .RW0_clk(mem_0_2_0_RW0_clk),
    .RW0_wdata(mem_0_2_0_RW0_wdata),
    .RW0_rdata(mem_0_2_0_RW0_rdata),
    .RW0_en(mem_0_2_0_RW0_en),
    .RW0_wmode(mem_0_2_0_RW0_wmode),
    .RW0_wmask(mem_0_2_0_RW0_wmask)
  );
  split_mem_ext mem_0_3_0 (
    .RW0_addr(mem_0_3_0_RW0_addr),
    .RW0_clk(mem_0_3_0_RW0_clk),
    .RW0_wdata(mem_0_3_0_RW0_wdata),
    .RW0_rdata(mem_0_3_0_RW0_rdata),
    .RW0_en(mem_0_3_0_RW0_en),
    .RW0_wmode(mem_0_3_0_RW0_wmode),
    .RW0_wmask(mem_0_3_0_RW0_wmask)
  );
  split_mem_ext mem_0_4_0 (
    .RW0_addr(mem_0_4_0_RW0_addr),
    .RW0_clk(mem_0_4_0_RW0_clk),
    .RW0_wdata(mem_0_4_0_RW0_wdata),
    .RW0_rdata(mem_0_4_0_RW0_rdata),
    .RW0_en(mem_0_4_0_RW0_en),
    .RW0_wmode(mem_0_4_0_RW0_wmode),
    .RW0_wmask(mem_0_4_0_RW0_wmask)
  );
  split_mem_ext mem_0_5_0 (
    .RW0_addr(mem_0_5_0_RW0_addr),
    .RW0_clk(mem_0_5_0_RW0_clk),
    .RW0_wdata(mem_0_5_0_RW0_wdata),
    .RW0_rdata(mem_0_5_0_RW0_rdata),
    .RW0_en(mem_0_5_0_RW0_en),
    .RW0_wmode(mem_0_5_0_RW0_wmode),
    .RW0_wmask(mem_0_5_0_RW0_wmask)
  );
  split_mem_ext mem_0_6_0 (
    .RW0_addr(mem_0_6_0_RW0_addr),
    .RW0_clk(mem_0_6_0_RW0_clk),
    .RW0_wdata(mem_0_6_0_RW0_wdata),
    .RW0_rdata(mem_0_6_0_RW0_rdata),
    .RW0_en(mem_0_6_0_RW0_en),
    .RW0_wmode(mem_0_6_0_RW0_wmode),
    .RW0_wmask(mem_0_6_0_RW0_wmask)
  );
  split_mem_ext mem_0_7_0 (
    .RW0_addr(mem_0_7_0_RW0_addr),
    .RW0_clk(mem_0_7_0_RW0_clk),
    .RW0_wdata(mem_0_7_0_RW0_wdata),
    .RW0_rdata(mem_0_7_0_RW0_rdata),
    .RW0_en(mem_0_7_0_RW0_en),
    .RW0_wmode(mem_0_7_0_RW0_wmode),
    .RW0_wmask(mem_0_7_0_RW0_wmask)
  );
  assign RW0_rdata = {RW0_rdata_0_7_0,_GEN_5};
  assign mem_0_0_0_RW0_addr = RW0_addr;
  assign mem_0_0_0_RW0_clk = RW0_clk;
  assign mem_0_0_0_RW0_wdata = RW0_wdata[7:0];
  assign mem_0_0_0_RW0_en = RW0_en;
  assign mem_0_0_0_RW0_wmode = RW0_wmode;
  assign mem_0_0_0_RW0_wmask = RW0_wmask[0];
  assign mem_0_1_0_RW0_addr = RW0_addr;
  assign mem_0_1_0_RW0_clk = RW0_clk;
  assign mem_0_1_0_RW0_wdata = RW0_wdata[15:8];
  assign mem_0_1_0_RW0_en = RW0_en;
  assign mem_0_1_0_RW0_wmode = RW0_wmode;
  assign mem_0_1_0_RW0_wmask = RW0_wmask[1];
  assign mem_0_2_0_RW0_addr = RW0_addr;
  assign mem_0_2_0_RW0_clk = RW0_clk;
  assign mem_0_2_0_RW0_wdata = RW0_wdata[23:16];
  assign mem_0_2_0_RW0_en = RW0_en;
  assign mem_0_2_0_RW0_wmode = RW0_wmode;
  assign mem_0_2_0_RW0_wmask = RW0_wmask[2];
  assign mem_0_3_0_RW0_addr = RW0_addr;
  assign mem_0_3_0_RW0_clk = RW0_clk;
  assign mem_0_3_0_RW0_wdata = RW0_wdata[31:24];
  assign mem_0_3_0_RW0_en = RW0_en;
  assign mem_0_3_0_RW0_wmode = RW0_wmode;
  assign mem_0_3_0_RW0_wmask = RW0_wmask[3];
  assign mem_0_4_0_RW0_addr = RW0_addr;
  assign mem_0_4_0_RW0_clk = RW0_clk;
  assign mem_0_4_0_RW0_wdata = RW0_wdata[39:32];
  assign mem_0_4_0_RW0_en = RW0_en;
  assign mem_0_4_0_RW0_wmode = RW0_wmode;
  assign mem_0_4_0_RW0_wmask = RW0_wmask[4];
  assign mem_0_5_0_RW0_addr = RW0_addr;
  assign mem_0_5_0_RW0_clk = RW0_clk;
  assign mem_0_5_0_RW0_wdata = RW0_wdata[47:40];
  assign mem_0_5_0_RW0_en = RW0_en;
  assign mem_0_5_0_RW0_wmode = RW0_wmode;
  assign mem_0_5_0_RW0_wmask = RW0_wmask[5];
  assign mem_0_6_0_RW0_addr = RW0_addr;
  assign mem_0_6_0_RW0_clk = RW0_clk;
  assign mem_0_6_0_RW0_wdata = RW0_wdata[55:48];
  assign mem_0_6_0_RW0_en = RW0_en;
  assign mem_0_6_0_RW0_wmode = RW0_wmode;
  assign mem_0_6_0_RW0_wmask = RW0_wmask[6];
  assign mem_0_7_0_RW0_addr = RW0_addr;
  assign mem_0_7_0_RW0_clk = RW0_clk;
  assign mem_0_7_0_RW0_wdata = RW0_wdata[63:56];
  assign mem_0_7_0_RW0_en = RW0_en;
  assign mem_0_7_0_RW0_wmode = RW0_wmode;
  assign mem_0_7_0_RW0_wmask = RW0_wmask[7];
endmodule
module split_mem_ext(
  input  [8:0] RW0_addr,
  input        RW0_clk,
  input  [7:0] RW0_wdata,
  output [7:0] RW0_rdata,
  input        RW0_en,
  input        RW0_wmode,
  input        RW0_wmask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:511];
  wire  ram_RW_0_r_en;
  wire [8:0] ram_RW_0_r_addr;
  wire [7:0] ram_RW_0_r_data;
  wire [7:0] ram_RW_0_w_data;
  wire [8:0] ram_RW_0_w_addr;
  wire  ram_RW_0_w_mask;
  wire  ram_RW_0_w_en;
  reg  ram_RW_0_r_en_pipe_0;
  reg [8:0] ram_RW_0_r_addr_pipe_0;
  wire  _GEN_0 = ~RW0_wmode;
  wire  _GEN_1 = ~RW0_wmode;
  assign ram_RW_0_r_en = ram_RW_0_r_en_pipe_0;
  assign ram_RW_0_r_addr = ram_RW_0_r_addr_pipe_0;
  assign ram_RW_0_r_data = ram[ram_RW_0_r_addr];
  assign ram_RW_0_w_data = RW0_wdata;
  assign ram_RW_0_w_addr = RW0_addr;
  assign ram_RW_0_w_mask = RW0_wmask;
  assign ram_RW_0_w_en = RW0_en & RW0_wmode;
  assign RW0_rdata = ram_RW_0_r_data;
  always @(posedge RW0_clk) begin
    if (ram_RW_0_w_en & ram_RW_0_w_mask) begin
      ram[ram_RW_0_w_addr] <= ram_RW_0_w_data;
    end
    ram_RW_0_r_en_pipe_0 <= RW0_en & ~RW0_wmode;
    if (RW0_en & ~RW0_wmode) begin
      ram_RW_0_r_addr_pipe_0 <= RW0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_RW_0_r_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_RW_0_r_addr_pipe_0 = _RAND_2[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
