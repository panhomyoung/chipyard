# Created by MC2 : Version 2012.02.00.d on 2025/06/20, 22:46:55

#*********************************************************************************************************************/
# Software       : TSMC MEMORY COMPILER tsn28hpcpuhdspsram_2012.02.00.d.170a						*/
# Technology     : TSMC 28nm CMOS LOGIC High Performance Compact Mobile Computing Plus 1P10M HKMG CU_ELK 0.9V				*/
#  Memory Type    : TSMC 28nm High Performance Compact Mobile Computing Plus Ultra High Density Single Port SRAM with d127 bit cell HVT periphery */
# Library Name   : ts1n28hpcpuhdhvtb32x50m4swbso (user specify : TS1N28HPCPUHDHVTB32X50M4SWBSO)				*/
# Library Version: 170a												*/
# Generated Time : 2025/06/20, 22:46:44										*/
#*********************************************************************************************************************/
#															*/
# STATEMENT OF USE													*/
#															*/
# This information contains confidential and proprietary information of TSMC.					*/
# No part of this information may be reproduced, transmitted, transcribed,						*/
# stored in a retrieval system, or translated into any human or computer						*/
# language, in any form or by any means, electronic, mechanical, magnetic,						*/
# optical, chemical, manual, or otherwise, without the prior written permission					*/
# of TSMC. This information was prepared for informational purpose and is for					*/
# use by TSMC's customers only. TSMC reserves the right to make changes in the					*/
# information at any time and without notice.									*/
#															*/
#*********************************************************************************************************************/
VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO TS1N28HPCPUHDHVTB32X50M4SWBSO
	CLASS BLOCK ;
	FOREIGN TS1N28HPCPUHDHVTB32X50M4SWBSO 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 18.890 BY 137.670 ;
	SYMMETRY X Y ;
	PIN AM[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 61.110 18.890 61.260 ;
			LAYER M3 ;
			RECT 18.710 61.110 18.890 61.260 ;
			LAYER M2 ;
			RECT 18.710 61.110 18.890 61.260 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.096800 LAYER M2 ;
		ANTENNAMAXAREACAR 5.155600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.755600 LAYER M3 ;
	END AM[0]

	PIN AM[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 62.100 18.890 62.250 ;
			LAYER M3 ;
			RECT 18.710 62.100 18.890 62.250 ;
			LAYER M1 ;
			RECT 18.710 62.100 18.890 62.250 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.096800 LAYER M2 ;
		ANTENNAMAXAREACAR 5.155600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.755600 LAYER M3 ;
	END AM[1]

	PIN AM[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 69.680 18.890 69.830 ;
			LAYER M3 ;
			RECT 18.710 69.680 18.890 69.830 ;
			LAYER M2 ;
			RECT 18.710 69.680 18.890 69.830 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.096800 LAYER M2 ;
		ANTENNAMAXAREACAR 5.155600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.755600 LAYER M3 ;
	END AM[2]

	PIN AM[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 70.320 18.890 70.470 ;
			LAYER M2 ;
			RECT 18.710 70.320 18.890 70.470 ;
			LAYER M1 ;
			RECT 18.710 70.320 18.890 70.470 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.096800 LAYER M2 ;
		ANTENNAMAXAREACAR 5.155600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.755600 LAYER M3 ;
	END AM[3]

	PIN AM[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 71.570 18.890 71.720 ;
			LAYER M1 ;
			RECT 18.710 71.570 18.890 71.720 ;
			LAYER M2 ;
			RECT 18.710 71.570 18.890 71.720 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.096800 LAYER M2 ;
		ANTENNAMAXAREACAR 5.155600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.755600 LAYER M3 ;
	END AM[4]

	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 61.440 18.890 61.590 ;
			LAYER M1 ;
			RECT 18.710 61.440 18.890 61.590 ;
			LAYER M3 ;
			RECT 18.710 61.440 18.890 61.590 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.670000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.123600 LAYER M2 ;
		ANTENNAMAXAREACAR 4.763600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.650000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.581800 LAYER M3 ;
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 61.770 18.890 61.920 ;
			LAYER M2 ;
			RECT 18.710 61.770 18.890 61.920 ;
			LAYER M1 ;
			RECT 18.710 61.770 18.890 61.920 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.670000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.123600 LAYER M2 ;
		ANTENNAMAXAREACAR 4.763600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.650000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.581800 LAYER M3 ;
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 69.220 18.890 69.370 ;
			LAYER M2 ;
			RECT 18.710 69.220 18.890 69.370 ;
			LAYER M1 ;
			RECT 18.710 69.220 18.890 69.370 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.670000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.123600 LAYER M2 ;
		ANTENNAMAXAREACAR 4.763600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.650000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.581800 LAYER M3 ;
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 70.780 18.890 70.930 ;
			LAYER M2 ;
			RECT 18.710 70.780 18.890 70.930 ;
			LAYER M3 ;
			RECT 18.710 70.780 18.890 70.930 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.670000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.123600 LAYER M2 ;
		ANTENNAMAXAREACAR 4.763600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.650000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.581800 LAYER M3 ;
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 71.110 18.890 71.260 ;
			LAYER M1 ;
			RECT 18.710 71.110 18.890 71.260 ;
			LAYER M2 ;
			RECT 18.710 71.110 18.890 71.260 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.670000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.433300 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.123600 LAYER M2 ;
		ANTENNAMAXAREACAR 4.763600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.650000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.581800 LAYER M3 ;
	END A[4]

	PIN BIST
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 74.065 18.890 74.215 ;
			LAYER M2 ;
			RECT 18.710 74.065 18.890 74.215 ;
			LAYER M1 ;
			RECT 18.710 74.065 18.890 74.215 ;
		END
		ANTENNAGATEAREA 0.120000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.115800 LAYER M1 ;
		ANTENNAMAXAREACAR 0.639600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.054200 LAYER VIA1 ;
		ANTENNAGATEAREA 0.120000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.091000 LAYER M2 ;
		ANTENNAMAXAREACAR 1.281200 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.108300 LAYER VIA2 ;
		ANTENNAGATEAREA 0.120000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.086400 LAYER M3 ;
		ANTENNAMAXAREACAR 1.506300 LAYER M3 ;
	END BIST

	PIN BWEBM[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 0.935 18.890 1.085 ;
			LAYER M3 ;
			RECT 18.710 0.935 18.890 1.085 ;
			LAYER M1 ;
			RECT 18.710 0.935 18.890 1.085 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[0]

	PIN BWEBM[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 24.135 18.890 24.285 ;
			LAYER M1 ;
			RECT 18.710 24.135 18.890 24.285 ;
			LAYER M2 ;
			RECT 18.710 24.135 18.890 24.285 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[10]

	PIN BWEBM[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 26.455 18.890 26.605 ;
			LAYER M1 ;
			RECT 18.710 26.455 18.890 26.605 ;
			LAYER M2 ;
			RECT 18.710 26.455 18.890 26.605 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[11]

	PIN BWEBM[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 28.775 18.890 28.925 ;
			LAYER M1 ;
			RECT 18.710 28.775 18.890 28.925 ;
			LAYER M3 ;
			RECT 18.710 28.775 18.890 28.925 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[12]

	PIN BWEBM[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 31.095 18.890 31.245 ;
			LAYER M3 ;
			RECT 18.710 31.095 18.890 31.245 ;
			LAYER M1 ;
			RECT 18.710 31.095 18.890 31.245 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[13]

	PIN BWEBM[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 33.415 18.890 33.565 ;
			LAYER M1 ;
			RECT 18.710 33.415 18.890 33.565 ;
			LAYER M2 ;
			RECT 18.710 33.415 18.890 33.565 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[14]

	PIN BWEBM[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 35.735 18.890 35.885 ;
			LAYER M2 ;
			RECT 18.710 35.735 18.890 35.885 ;
			LAYER M3 ;
			RECT 18.710 35.735 18.890 35.885 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[15]

	PIN BWEBM[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 38.055 18.890 38.205 ;
			LAYER M2 ;
			RECT 18.710 38.055 18.890 38.205 ;
			LAYER M1 ;
			RECT 18.710 38.055 18.890 38.205 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[16]

	PIN BWEBM[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 40.375 18.890 40.525 ;
			LAYER M2 ;
			RECT 18.710 40.375 18.890 40.525 ;
			LAYER M3 ;
			RECT 18.710 40.375 18.890 40.525 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[17]

	PIN BWEBM[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 42.695 18.890 42.845 ;
			LAYER M1 ;
			RECT 18.710 42.695 18.890 42.845 ;
			LAYER M3 ;
			RECT 18.710 42.695 18.890 42.845 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[18]

	PIN BWEBM[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 45.015 18.890 45.165 ;
			LAYER M2 ;
			RECT 18.710 45.015 18.890 45.165 ;
			LAYER M3 ;
			RECT 18.710 45.015 18.890 45.165 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[19]

	PIN BWEBM[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 3.255 18.890 3.405 ;
			LAYER M2 ;
			RECT 18.710 3.255 18.890 3.405 ;
			LAYER M3 ;
			RECT 18.710 3.255 18.890 3.405 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[1]

	PIN BWEBM[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 47.335 18.890 47.485 ;
			LAYER M1 ;
			RECT 18.710 47.335 18.890 47.485 ;
			LAYER M2 ;
			RECT 18.710 47.335 18.890 47.485 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[20]

	PIN BWEBM[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 49.655 18.890 49.805 ;
			LAYER M2 ;
			RECT 18.710 49.655 18.890 49.805 ;
			LAYER M3 ;
			RECT 18.710 49.655 18.890 49.805 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[21]

	PIN BWEBM[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 51.975 18.890 52.125 ;
			LAYER M3 ;
			RECT 18.710 51.975 18.890 52.125 ;
			LAYER M2 ;
			RECT 18.710 51.975 18.890 52.125 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[22]

	PIN BWEBM[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 54.295 18.890 54.445 ;
			LAYER M3 ;
			RECT 18.710 54.295 18.890 54.445 ;
			LAYER M1 ;
			RECT 18.710 54.295 18.890 54.445 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[23]

	PIN BWEBM[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 56.615 18.890 56.765 ;
			LAYER M1 ;
			RECT 18.710 56.615 18.890 56.765 ;
			LAYER M3 ;
			RECT 18.710 56.615 18.890 56.765 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[24]

	PIN BWEBM[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 78.935 18.890 79.085 ;
			LAYER M1 ;
			RECT 18.710 78.935 18.890 79.085 ;
			LAYER M2 ;
			RECT 18.710 78.935 18.890 79.085 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[25]

	PIN BWEBM[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 81.255 18.890 81.405 ;
			LAYER M2 ;
			RECT 18.710 81.255 18.890 81.405 ;
			LAYER M3 ;
			RECT 18.710 81.255 18.890 81.405 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[26]

	PIN BWEBM[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 83.575 18.890 83.725 ;
			LAYER M1 ;
			RECT 18.710 83.575 18.890 83.725 ;
			LAYER M2 ;
			RECT 18.710 83.575 18.890 83.725 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[27]

	PIN BWEBM[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 85.895 18.890 86.045 ;
			LAYER M3 ;
			RECT 18.710 85.895 18.890 86.045 ;
			LAYER M1 ;
			RECT 18.710 85.895 18.890 86.045 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[28]

	PIN BWEBM[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 88.215 18.890 88.365 ;
			LAYER M3 ;
			RECT 18.710 88.215 18.890 88.365 ;
			LAYER M1 ;
			RECT 18.710 88.215 18.890 88.365 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[29]

	PIN BWEBM[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 5.575 18.890 5.725 ;
			LAYER M3 ;
			RECT 18.710 5.575 18.890 5.725 ;
			LAYER M2 ;
			RECT 18.710 5.575 18.890 5.725 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[2]

	PIN BWEBM[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 90.535 18.890 90.685 ;
			LAYER M1 ;
			RECT 18.710 90.535 18.890 90.685 ;
			LAYER M2 ;
			RECT 18.710 90.535 18.890 90.685 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[30]

	PIN BWEBM[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 92.855 18.890 93.005 ;
			LAYER M1 ;
			RECT 18.710 92.855 18.890 93.005 ;
			LAYER M2 ;
			RECT 18.710 92.855 18.890 93.005 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[31]

	PIN BWEBM[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 95.175 18.890 95.325 ;
			LAYER M2 ;
			RECT 18.710 95.175 18.890 95.325 ;
			LAYER M3 ;
			RECT 18.710 95.175 18.890 95.325 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[32]

	PIN BWEBM[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 97.495 18.890 97.645 ;
			LAYER M2 ;
			RECT 18.710 97.495 18.890 97.645 ;
			LAYER M3 ;
			RECT 18.710 97.495 18.890 97.645 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[33]

	PIN BWEBM[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 99.815 18.890 99.965 ;
			LAYER M1 ;
			RECT 18.710 99.815 18.890 99.965 ;
			LAYER M2 ;
			RECT 18.710 99.815 18.890 99.965 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[34]

	PIN BWEBM[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 102.135 18.890 102.285 ;
			LAYER M2 ;
			RECT 18.710 102.135 18.890 102.285 ;
			LAYER M1 ;
			RECT 18.710 102.135 18.890 102.285 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[35]

	PIN BWEBM[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 104.455 18.890 104.605 ;
			LAYER M2 ;
			RECT 18.710 104.455 18.890 104.605 ;
			LAYER M1 ;
			RECT 18.710 104.455 18.890 104.605 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[36]

	PIN BWEBM[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 106.775 18.890 106.925 ;
			LAYER M2 ;
			RECT 18.710 106.775 18.890 106.925 ;
			LAYER M3 ;
			RECT 18.710 106.775 18.890 106.925 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[37]

	PIN BWEBM[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 109.095 18.890 109.245 ;
			LAYER M2 ;
			RECT 18.710 109.095 18.890 109.245 ;
			LAYER M3 ;
			RECT 18.710 109.095 18.890 109.245 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[38]

	PIN BWEBM[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 111.415 18.890 111.565 ;
			LAYER M2 ;
			RECT 18.710 111.415 18.890 111.565 ;
			LAYER M3 ;
			RECT 18.710 111.415 18.890 111.565 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[39]

	PIN BWEBM[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 7.895 18.890 8.045 ;
			LAYER M2 ;
			RECT 18.710 7.895 18.890 8.045 ;
			LAYER M3 ;
			RECT 18.710 7.895 18.890 8.045 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[3]

	PIN BWEBM[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 113.735 18.890 113.885 ;
			LAYER M3 ;
			RECT 18.710 113.735 18.890 113.885 ;
			LAYER M2 ;
			RECT 18.710 113.735 18.890 113.885 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[40]

	PIN BWEBM[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 116.055 18.890 116.205 ;
			LAYER M3 ;
			RECT 18.710 116.055 18.890 116.205 ;
			LAYER M1 ;
			RECT 18.710 116.055 18.890 116.205 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[41]

	PIN BWEBM[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 118.375 18.890 118.525 ;
			LAYER M3 ;
			RECT 18.710 118.375 18.890 118.525 ;
			LAYER M1 ;
			RECT 18.710 118.375 18.890 118.525 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[42]

	PIN BWEBM[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 120.695 18.890 120.845 ;
			LAYER M2 ;
			RECT 18.710 120.695 18.890 120.845 ;
			LAYER M1 ;
			RECT 18.710 120.695 18.890 120.845 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[43]

	PIN BWEBM[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 123.015 18.890 123.165 ;
			LAYER M2 ;
			RECT 18.710 123.015 18.890 123.165 ;
			LAYER M1 ;
			RECT 18.710 123.015 18.890 123.165 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[44]

	PIN BWEBM[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 125.335 18.890 125.485 ;
			LAYER M3 ;
			RECT 18.710 125.335 18.890 125.485 ;
			LAYER M2 ;
			RECT 18.710 125.335 18.890 125.485 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[45]

	PIN BWEBM[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 127.655 18.890 127.805 ;
			LAYER M1 ;
			RECT 18.710 127.655 18.890 127.805 ;
			LAYER M2 ;
			RECT 18.710 127.655 18.890 127.805 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[46]

	PIN BWEBM[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 129.975 18.890 130.125 ;
			LAYER M1 ;
			RECT 18.710 129.975 18.890 130.125 ;
			LAYER M3 ;
			RECT 18.710 129.975 18.890 130.125 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[47]

	PIN BWEBM[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 132.295 18.890 132.445 ;
			LAYER M3 ;
			RECT 18.710 132.295 18.890 132.445 ;
			LAYER M1 ;
			RECT 18.710 132.295 18.890 132.445 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[48]

	PIN BWEBM[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 134.615 18.890 134.765 ;
			LAYER M3 ;
			RECT 18.710 134.615 18.890 134.765 ;
			LAYER M2 ;
			RECT 18.710 134.615 18.890 134.765 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[49]

	PIN BWEBM[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 10.215 18.890 10.365 ;
			LAYER M3 ;
			RECT 18.710 10.215 18.890 10.365 ;
			LAYER M1 ;
			RECT 18.710 10.215 18.890 10.365 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[4]

	PIN BWEBM[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 12.535 18.890 12.685 ;
			LAYER M1 ;
			RECT 18.710 12.535 18.890 12.685 ;
			LAYER M3 ;
			RECT 18.710 12.535 18.890 12.685 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[5]

	PIN BWEBM[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 14.855 18.890 15.005 ;
			LAYER M2 ;
			RECT 18.710 14.855 18.890 15.005 ;
			LAYER M1 ;
			RECT 18.710 14.855 18.890 15.005 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[6]

	PIN BWEBM[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 17.175 18.890 17.325 ;
			LAYER M2 ;
			RECT 18.710 17.175 18.890 17.325 ;
			LAYER M3 ;
			RECT 18.710 17.175 18.890 17.325 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[7]

	PIN BWEBM[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 19.495 18.890 19.645 ;
			LAYER M2 ;
			RECT 18.710 19.495 18.890 19.645 ;
			LAYER M1 ;
			RECT 18.710 19.495 18.890 19.645 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[8]

	PIN BWEBM[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 21.815 18.890 21.965 ;
			LAYER M3 ;
			RECT 18.710 21.815 18.890 21.965 ;
			LAYER M2 ;
			RECT 18.710 21.815 18.890 21.965 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 12.682300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 13.067700 LAYER M3 ;
	END BWEBM[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 1.265 18.890 1.415 ;
			LAYER M1 ;
			RECT 18.710 1.265 18.890 1.415 ;
			LAYER M2 ;
			RECT 18.710 1.265 18.890 1.415 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[0]

	PIN BWEB[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 24.465 18.890 24.615 ;
			LAYER M1 ;
			RECT 18.710 24.465 18.890 24.615 ;
			LAYER M3 ;
			RECT 18.710 24.465 18.890 24.615 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[10]

	PIN BWEB[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 26.785 18.890 26.935 ;
			LAYER M2 ;
			RECT 18.710 26.785 18.890 26.935 ;
			LAYER M3 ;
			RECT 18.710 26.785 18.890 26.935 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[11]

	PIN BWEB[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 29.105 18.890 29.255 ;
			LAYER M1 ;
			RECT 18.710 29.105 18.890 29.255 ;
			LAYER M3 ;
			RECT 18.710 29.105 18.890 29.255 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[12]

	PIN BWEB[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 31.425 18.890 31.575 ;
			LAYER M2 ;
			RECT 18.710 31.425 18.890 31.575 ;
			LAYER M1 ;
			RECT 18.710 31.425 18.890 31.575 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[13]

	PIN BWEB[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 33.745 18.890 33.895 ;
			LAYER M3 ;
			RECT 18.710 33.745 18.890 33.895 ;
			LAYER M2 ;
			RECT 18.710 33.745 18.890 33.895 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[14]

	PIN BWEB[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 36.065 18.890 36.215 ;
			LAYER M1 ;
			RECT 18.710 36.065 18.890 36.215 ;
			LAYER M2 ;
			RECT 18.710 36.065 18.890 36.215 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[15]

	PIN BWEB[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 38.385 18.890 38.535 ;
			LAYER M2 ;
			RECT 18.710 38.385 18.890 38.535 ;
			LAYER M3 ;
			RECT 18.710 38.385 18.890 38.535 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[16]

	PIN BWEB[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 40.705 18.890 40.855 ;
			LAYER M3 ;
			RECT 18.710 40.705 18.890 40.855 ;
			LAYER M1 ;
			RECT 18.710 40.705 18.890 40.855 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[17]

	PIN BWEB[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 43.025 18.890 43.175 ;
			LAYER M2 ;
			RECT 18.710 43.025 18.890 43.175 ;
			LAYER M3 ;
			RECT 18.710 43.025 18.890 43.175 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[18]

	PIN BWEB[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 45.345 18.890 45.495 ;
			LAYER M1 ;
			RECT 18.710 45.345 18.890 45.495 ;
			LAYER M3 ;
			RECT 18.710 45.345 18.890 45.495 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[19]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 3.585 18.890 3.735 ;
			LAYER M1 ;
			RECT 18.710 3.585 18.890 3.735 ;
			LAYER M3 ;
			RECT 18.710 3.585 18.890 3.735 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[1]

	PIN BWEB[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 47.665 18.890 47.815 ;
			LAYER M3 ;
			RECT 18.710 47.665 18.890 47.815 ;
			LAYER M1 ;
			RECT 18.710 47.665 18.890 47.815 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[20]

	PIN BWEB[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 49.985 18.890 50.135 ;
			LAYER M2 ;
			RECT 18.710 49.985 18.890 50.135 ;
			LAYER M3 ;
			RECT 18.710 49.985 18.890 50.135 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[21]

	PIN BWEB[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 52.305 18.890 52.455 ;
			LAYER M1 ;
			RECT 18.710 52.305 18.890 52.455 ;
			LAYER M3 ;
			RECT 18.710 52.305 18.890 52.455 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[22]

	PIN BWEB[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 54.625 18.890 54.775 ;
			LAYER M2 ;
			RECT 18.710 54.625 18.890 54.775 ;
			LAYER M1 ;
			RECT 18.710 54.625 18.890 54.775 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[23]

	PIN BWEB[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 56.945 18.890 57.095 ;
			LAYER M3 ;
			RECT 18.710 56.945 18.890 57.095 ;
			LAYER M2 ;
			RECT 18.710 56.945 18.890 57.095 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[24]

	PIN BWEB[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 79.265 18.890 79.415 ;
			LAYER M1 ;
			RECT 18.710 79.265 18.890 79.415 ;
			LAYER M3 ;
			RECT 18.710 79.265 18.890 79.415 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[25]

	PIN BWEB[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 81.585 18.890 81.735 ;
			LAYER M1 ;
			RECT 18.710 81.585 18.890 81.735 ;
			LAYER M2 ;
			RECT 18.710 81.585 18.890 81.735 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[26]

	PIN BWEB[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 83.905 18.890 84.055 ;
			LAYER M2 ;
			RECT 18.710 83.905 18.890 84.055 ;
			LAYER M1 ;
			RECT 18.710 83.905 18.890 84.055 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[27]

	PIN BWEB[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 86.225 18.890 86.375 ;
			LAYER M2 ;
			RECT 18.710 86.225 18.890 86.375 ;
			LAYER M3 ;
			RECT 18.710 86.225 18.890 86.375 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[28]

	PIN BWEB[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 88.545 18.890 88.695 ;
			LAYER M2 ;
			RECT 18.710 88.545 18.890 88.695 ;
			LAYER M3 ;
			RECT 18.710 88.545 18.890 88.695 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[29]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 5.905 18.890 6.055 ;
			LAYER M3 ;
			RECT 18.710 5.905 18.890 6.055 ;
			LAYER M1 ;
			RECT 18.710 5.905 18.890 6.055 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[2]

	PIN BWEB[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 90.865 18.890 91.015 ;
			LAYER M1 ;
			RECT 18.710 90.865 18.890 91.015 ;
			LAYER M3 ;
			RECT 18.710 90.865 18.890 91.015 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[30]

	PIN BWEB[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 93.185 18.890 93.335 ;
			LAYER M1 ;
			RECT 18.710 93.185 18.890 93.335 ;
			LAYER M2 ;
			RECT 18.710 93.185 18.890 93.335 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[31]

	PIN BWEB[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 95.505 18.890 95.655 ;
			LAYER M2 ;
			RECT 18.710 95.505 18.890 95.655 ;
			LAYER M3 ;
			RECT 18.710 95.505 18.890 95.655 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[32]

	PIN BWEB[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 97.825 18.890 97.975 ;
			LAYER M3 ;
			RECT 18.710 97.825 18.890 97.975 ;
			LAYER M1 ;
			RECT 18.710 97.825 18.890 97.975 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[33]

	PIN BWEB[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 100.145 18.890 100.295 ;
			LAYER M2 ;
			RECT 18.710 100.145 18.890 100.295 ;
			LAYER M1 ;
			RECT 18.710 100.145 18.890 100.295 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[34]

	PIN BWEB[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 102.465 18.890 102.615 ;
			LAYER M3 ;
			RECT 18.710 102.465 18.890 102.615 ;
			LAYER M2 ;
			RECT 18.710 102.465 18.890 102.615 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[35]

	PIN BWEB[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 104.785 18.890 104.935 ;
			LAYER M2 ;
			RECT 18.710 104.785 18.890 104.935 ;
			LAYER M3 ;
			RECT 18.710 104.785 18.890 104.935 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[36]

	PIN BWEB[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 107.105 18.890 107.255 ;
			LAYER M1 ;
			RECT 18.710 107.105 18.890 107.255 ;
			LAYER M2 ;
			RECT 18.710 107.105 18.890 107.255 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[37]

	PIN BWEB[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 109.425 18.890 109.575 ;
			LAYER M3 ;
			RECT 18.710 109.425 18.890 109.575 ;
			LAYER M2 ;
			RECT 18.710 109.425 18.890 109.575 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[38]

	PIN BWEB[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 111.745 18.890 111.895 ;
			LAYER M2 ;
			RECT 18.710 111.745 18.890 111.895 ;
			LAYER M3 ;
			RECT 18.710 111.745 18.890 111.895 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[39]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 8.225 18.890 8.375 ;
			LAYER M2 ;
			RECT 18.710 8.225 18.890 8.375 ;
			LAYER M3 ;
			RECT 18.710 8.225 18.890 8.375 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[3]

	PIN BWEB[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 114.065 18.890 114.215 ;
			LAYER M1 ;
			RECT 18.710 114.065 18.890 114.215 ;
			LAYER M2 ;
			RECT 18.710 114.065 18.890 114.215 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[40]

	PIN BWEB[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 116.385 18.890 116.535 ;
			LAYER M1 ;
			RECT 18.710 116.385 18.890 116.535 ;
			LAYER M2 ;
			RECT 18.710 116.385 18.890 116.535 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[41]

	PIN BWEB[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 118.705 18.890 118.855 ;
			LAYER M2 ;
			RECT 18.710 118.705 18.890 118.855 ;
			LAYER M3 ;
			RECT 18.710 118.705 18.890 118.855 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[42]

	PIN BWEB[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 121.025 18.890 121.175 ;
			LAYER M1 ;
			RECT 18.710 121.025 18.890 121.175 ;
			LAYER M2 ;
			RECT 18.710 121.025 18.890 121.175 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[43]

	PIN BWEB[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 123.345 18.890 123.495 ;
			LAYER M3 ;
			RECT 18.710 123.345 18.890 123.495 ;
			LAYER M1 ;
			RECT 18.710 123.345 18.890 123.495 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[44]

	PIN BWEB[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 125.665 18.890 125.815 ;
			LAYER M2 ;
			RECT 18.710 125.665 18.890 125.815 ;
			LAYER M3 ;
			RECT 18.710 125.665 18.890 125.815 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[45]

	PIN BWEB[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 127.985 18.890 128.135 ;
			LAYER M3 ;
			RECT 18.710 127.985 18.890 128.135 ;
			LAYER M1 ;
			RECT 18.710 127.985 18.890 128.135 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[46]

	PIN BWEB[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 130.305 18.890 130.455 ;
			LAYER M2 ;
			RECT 18.710 130.305 18.890 130.455 ;
			LAYER M1 ;
			RECT 18.710 130.305 18.890 130.455 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[47]

	PIN BWEB[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 132.625 18.890 132.775 ;
			LAYER M2 ;
			RECT 18.710 132.625 18.890 132.775 ;
			LAYER M1 ;
			RECT 18.710 132.625 18.890 132.775 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[48]

	PIN BWEB[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 134.945 18.890 135.095 ;
			LAYER M3 ;
			RECT 18.710 134.945 18.890 135.095 ;
			LAYER M1 ;
			RECT 18.710 134.945 18.890 135.095 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[49]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 10.545 18.890 10.695 ;
			LAYER M1 ;
			RECT 18.710 10.545 18.890 10.695 ;
			LAYER M2 ;
			RECT 18.710 10.545 18.890 10.695 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 12.865 18.890 13.015 ;
			LAYER M2 ;
			RECT 18.710 12.865 18.890 13.015 ;
			LAYER M1 ;
			RECT 18.710 12.865 18.890 13.015 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 15.185 18.890 15.335 ;
			LAYER M2 ;
			RECT 18.710 15.185 18.890 15.335 ;
			LAYER M1 ;
			RECT 18.710 15.185 18.890 15.335 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 17.505 18.890 17.655 ;
			LAYER M2 ;
			RECT 18.710 17.505 18.890 17.655 ;
			LAYER M3 ;
			RECT 18.710 17.505 18.890 17.655 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[7]

	PIN BWEB[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 19.825 18.890 19.975 ;
			LAYER M2 ;
			RECT 18.710 19.825 18.890 19.975 ;
			LAYER M3 ;
			RECT 18.710 19.825 18.890 19.975 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[8]

	PIN BWEB[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 22.145 18.890 22.295 ;
			LAYER M1 ;
			RECT 18.710 22.145 18.890 22.295 ;
			LAYER M3 ;
			RECT 18.710 22.145 18.890 22.295 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.086200 LAYER M1 ;
		ANTENNAMAXAREACAR 8.984400 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118700 LAYER M2 ;
		ANTENNAMAXAREACAR 11.796900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.052200 LAYER M3 ;
		ANTENNAMAXAREACAR 16.010400 LAYER M3 ;
	END BWEB[9]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 72.670 18.890 72.820 ;
			LAYER M3 ;
			RECT 18.710 72.670 18.890 72.820 ;
			LAYER M2 ;
			RECT 18.710 72.670 18.890 72.820 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.670000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.393900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.118200 LAYER M2 ;
		ANTENNAMAXAREACAR 4.503000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.590900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.321200 LAYER M3 ;
	END CEB

	PIN CEBM
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 72.210 18.890 72.360 ;
			LAYER M3 ;
			RECT 18.710 72.210 18.890 72.360 ;
			LAYER M2 ;
			RECT 18.710 72.210 18.890 72.360 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.092700 LAYER M2 ;
		ANTENNAMAXAREACAR 5.066700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.666700 LAYER M3 ;
	END CEBM

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 76.070 18.890 76.220 ;
			LAYER M1 ;
			RECT 18.710 76.070 18.890 76.220 ;
			LAYER M3 ;
			RECT 18.710 76.070 18.890 76.220 ;
		END
		ANTENNAGATEAREA 0.149100 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.229300 LAYER M1 ;
		ANTENNAMAXAREACAR 1.425900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.045500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.408800 LAYER VIA1 ;
		ANTENNAGATEAREA 0.149100 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.059500 LAYER M2 ;
		ANTENNAMAXAREACAR 8.761900 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.642000 LAYER VIA2 ;
		ANTENNAGATEAREA 0.149100 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.113500 LAYER M3 ;
		ANTENNAMAXAREACAR 9.523100 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 0.496000 LAYER VIA3 ;
		ANTENNAGATEAREA 0.149100 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 12.551900 LAYER M4 ;
		ANTENNAMAXAREACAR 88.259300 LAYER M4 ;
	END CLK

	PIN DM[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 2.905 18.890 3.055 ;
			LAYER M3 ;
			RECT 18.710 2.905 18.890 3.055 ;
			LAYER M1 ;
			RECT 18.710 2.905 18.890 3.055 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[0]

	PIN DM[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 26.105 18.890 26.255 ;
			LAYER M2 ;
			RECT 18.710 26.105 18.890 26.255 ;
			LAYER M1 ;
			RECT 18.710 26.105 18.890 26.255 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[10]

	PIN DM[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 28.425 18.890 28.575 ;
			LAYER M2 ;
			RECT 18.710 28.425 18.890 28.575 ;
			LAYER M1 ;
			RECT 18.710 28.425 18.890 28.575 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[11]

	PIN DM[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 30.745 18.890 30.895 ;
			LAYER M1 ;
			RECT 18.710 30.745 18.890 30.895 ;
			LAYER M2 ;
			RECT 18.710 30.745 18.890 30.895 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[12]

	PIN DM[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 33.065 18.890 33.215 ;
			LAYER M2 ;
			RECT 18.710 33.065 18.890 33.215 ;
			LAYER M1 ;
			RECT 18.710 33.065 18.890 33.215 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[13]

	PIN DM[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 35.385 18.890 35.535 ;
			LAYER M1 ;
			RECT 18.710 35.385 18.890 35.535 ;
			LAYER M2 ;
			RECT 18.710 35.385 18.890 35.535 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[14]

	PIN DM[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 37.705 18.890 37.855 ;
			LAYER M3 ;
			RECT 18.710 37.705 18.890 37.855 ;
			LAYER M2 ;
			RECT 18.710 37.705 18.890 37.855 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[15]

	PIN DM[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 40.025 18.890 40.175 ;
			LAYER M2 ;
			RECT 18.710 40.025 18.890 40.175 ;
			LAYER M1 ;
			RECT 18.710 40.025 18.890 40.175 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[16]

	PIN DM[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 42.345 18.890 42.495 ;
			LAYER M3 ;
			RECT 18.710 42.345 18.890 42.495 ;
			LAYER M1 ;
			RECT 18.710 42.345 18.890 42.495 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[17]

	PIN DM[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 44.665 18.890 44.815 ;
			LAYER M3 ;
			RECT 18.710 44.665 18.890 44.815 ;
			LAYER M2 ;
			RECT 18.710 44.665 18.890 44.815 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[18]

	PIN DM[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 46.985 18.890 47.135 ;
			LAYER M2 ;
			RECT 18.710 46.985 18.890 47.135 ;
			LAYER M1 ;
			RECT 18.710 46.985 18.890 47.135 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[19]

	PIN DM[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 5.225 18.890 5.375 ;
			LAYER M2 ;
			RECT 18.710 5.225 18.890 5.375 ;
			LAYER M1 ;
			RECT 18.710 5.225 18.890 5.375 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[1]

	PIN DM[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 49.305 18.890 49.455 ;
			LAYER M3 ;
			RECT 18.710 49.305 18.890 49.455 ;
			LAYER M2 ;
			RECT 18.710 49.305 18.890 49.455 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[20]

	PIN DM[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 51.625 18.890 51.775 ;
			LAYER M1 ;
			RECT 18.710 51.625 18.890 51.775 ;
			LAYER M3 ;
			RECT 18.710 51.625 18.890 51.775 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[21]

	PIN DM[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 53.945 18.890 54.095 ;
			LAYER M2 ;
			RECT 18.710 53.945 18.890 54.095 ;
			LAYER M1 ;
			RECT 18.710 53.945 18.890 54.095 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[22]

	PIN DM[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 56.265 18.890 56.415 ;
			LAYER M1 ;
			RECT 18.710 56.265 18.890 56.415 ;
			LAYER M2 ;
			RECT 18.710 56.265 18.890 56.415 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[23]

	PIN DM[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 58.585 18.890 58.735 ;
			LAYER M1 ;
			RECT 18.710 58.585 18.890 58.735 ;
			LAYER M2 ;
			RECT 18.710 58.585 18.890 58.735 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[24]

	PIN DM[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 80.905 18.890 81.055 ;
			LAYER M1 ;
			RECT 18.710 80.905 18.890 81.055 ;
			LAYER M2 ;
			RECT 18.710 80.905 18.890 81.055 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[25]

	PIN DM[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 83.225 18.890 83.375 ;
			LAYER M2 ;
			RECT 18.710 83.225 18.890 83.375 ;
			LAYER M3 ;
			RECT 18.710 83.225 18.890 83.375 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[26]

	PIN DM[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 85.545 18.890 85.695 ;
			LAYER M3 ;
			RECT 18.710 85.545 18.890 85.695 ;
			LAYER M2 ;
			RECT 18.710 85.545 18.890 85.695 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[27]

	PIN DM[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 87.865 18.890 88.015 ;
			LAYER M2 ;
			RECT 18.710 87.865 18.890 88.015 ;
			LAYER M3 ;
			RECT 18.710 87.865 18.890 88.015 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[28]

	PIN DM[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 90.185 18.890 90.335 ;
			LAYER M2 ;
			RECT 18.710 90.185 18.890 90.335 ;
			LAYER M1 ;
			RECT 18.710 90.185 18.890 90.335 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[29]

	PIN DM[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 7.545 18.890 7.695 ;
			LAYER M2 ;
			RECT 18.710 7.545 18.890 7.695 ;
			LAYER M3 ;
			RECT 18.710 7.545 18.890 7.695 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[2]

	PIN DM[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 92.505 18.890 92.655 ;
			LAYER M3 ;
			RECT 18.710 92.505 18.890 92.655 ;
			LAYER M1 ;
			RECT 18.710 92.505 18.890 92.655 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[30]

	PIN DM[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 94.825 18.890 94.975 ;
			LAYER M2 ;
			RECT 18.710 94.825 18.890 94.975 ;
			LAYER M3 ;
			RECT 18.710 94.825 18.890 94.975 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[31]

	PIN DM[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 97.145 18.890 97.295 ;
			LAYER M2 ;
			RECT 18.710 97.145 18.890 97.295 ;
			LAYER M1 ;
			RECT 18.710 97.145 18.890 97.295 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[32]

	PIN DM[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 99.465 18.890 99.615 ;
			LAYER M1 ;
			RECT 18.710 99.465 18.890 99.615 ;
			LAYER M3 ;
			RECT 18.710 99.465 18.890 99.615 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[33]

	PIN DM[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 101.785 18.890 101.935 ;
			LAYER M1 ;
			RECT 18.710 101.785 18.890 101.935 ;
			LAYER M3 ;
			RECT 18.710 101.785 18.890 101.935 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[34]

	PIN DM[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 104.105 18.890 104.255 ;
			LAYER M1 ;
			RECT 18.710 104.105 18.890 104.255 ;
			LAYER M3 ;
			RECT 18.710 104.105 18.890 104.255 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[35]

	PIN DM[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 106.425 18.890 106.575 ;
			LAYER M1 ;
			RECT 18.710 106.425 18.890 106.575 ;
			LAYER M2 ;
			RECT 18.710 106.425 18.890 106.575 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[36]

	PIN DM[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 108.745 18.890 108.895 ;
			LAYER M1 ;
			RECT 18.710 108.745 18.890 108.895 ;
			LAYER M3 ;
			RECT 18.710 108.745 18.890 108.895 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[37]

	PIN DM[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 111.065 18.890 111.215 ;
			LAYER M2 ;
			RECT 18.710 111.065 18.890 111.215 ;
			LAYER M1 ;
			RECT 18.710 111.065 18.890 111.215 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[38]

	PIN DM[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 113.385 18.890 113.535 ;
			LAYER M3 ;
			RECT 18.710 113.385 18.890 113.535 ;
			LAYER M2 ;
			RECT 18.710 113.385 18.890 113.535 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[39]

	PIN DM[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 9.865 18.890 10.015 ;
			LAYER M1 ;
			RECT 18.710 9.865 18.890 10.015 ;
			LAYER M2 ;
			RECT 18.710 9.865 18.890 10.015 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[3]

	PIN DM[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 115.705 18.890 115.855 ;
			LAYER M2 ;
			RECT 18.710 115.705 18.890 115.855 ;
			LAYER M1 ;
			RECT 18.710 115.705 18.890 115.855 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[40]

	PIN DM[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 118.025 18.890 118.175 ;
			LAYER M2 ;
			RECT 18.710 118.025 18.890 118.175 ;
			LAYER M1 ;
			RECT 18.710 118.025 18.890 118.175 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[41]

	PIN DM[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 120.345 18.890 120.495 ;
			LAYER M3 ;
			RECT 18.710 120.345 18.890 120.495 ;
			LAYER M2 ;
			RECT 18.710 120.345 18.890 120.495 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[42]

	PIN DM[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 122.665 18.890 122.815 ;
			LAYER M1 ;
			RECT 18.710 122.665 18.890 122.815 ;
			LAYER M3 ;
			RECT 18.710 122.665 18.890 122.815 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[43]

	PIN DM[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 124.985 18.890 125.135 ;
			LAYER M2 ;
			RECT 18.710 124.985 18.890 125.135 ;
			LAYER M3 ;
			RECT 18.710 124.985 18.890 125.135 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[44]

	PIN DM[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 127.305 18.890 127.455 ;
			LAYER M3 ;
			RECT 18.710 127.305 18.890 127.455 ;
			LAYER M2 ;
			RECT 18.710 127.305 18.890 127.455 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[45]

	PIN DM[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 129.625 18.890 129.775 ;
			LAYER M3 ;
			RECT 18.710 129.625 18.890 129.775 ;
			LAYER M1 ;
			RECT 18.710 129.625 18.890 129.775 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[46]

	PIN DM[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 131.945 18.890 132.095 ;
			LAYER M1 ;
			RECT 18.710 131.945 18.890 132.095 ;
			LAYER M2 ;
			RECT 18.710 131.945 18.890 132.095 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[47]

	PIN DM[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 134.265 18.890 134.415 ;
			LAYER M2 ;
			RECT 18.710 134.265 18.890 134.415 ;
			LAYER M1 ;
			RECT 18.710 134.265 18.890 134.415 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[48]

	PIN DM[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 136.585 18.890 136.735 ;
			LAYER M2 ;
			RECT 18.710 136.585 18.890 136.735 ;
			LAYER M1 ;
			RECT 18.710 136.585 18.890 136.735 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[49]

	PIN DM[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 12.185 18.890 12.335 ;
			LAYER M2 ;
			RECT 18.710 12.185 18.890 12.335 ;
			LAYER M3 ;
			RECT 18.710 12.185 18.890 12.335 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[4]

	PIN DM[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 14.505 18.890 14.655 ;
			LAYER M3 ;
			RECT 18.710 14.505 18.890 14.655 ;
			LAYER M2 ;
			RECT 18.710 14.505 18.890 14.655 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[5]

	PIN DM[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 16.825 18.890 16.975 ;
			LAYER M1 ;
			RECT 18.710 16.825 18.890 16.975 ;
			LAYER M3 ;
			RECT 18.710 16.825 18.890 16.975 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[6]

	PIN DM[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 19.145 18.890 19.295 ;
			LAYER M1 ;
			RECT 18.710 19.145 18.890 19.295 ;
			LAYER M3 ;
			RECT 18.710 19.145 18.890 19.295 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[7]

	PIN DM[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 21.465 18.890 21.615 ;
			LAYER M1 ;
			RECT 18.710 21.465 18.890 21.615 ;
			LAYER M2 ;
			RECT 18.710 21.465 18.890 21.615 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[8]

	PIN DM[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 23.785 18.890 23.935 ;
			LAYER M2 ;
			RECT 18.710 23.785 18.890 23.935 ;
			LAYER M1 ;
			RECT 18.710 23.785 18.890 23.935 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.080900 LAYER M1 ;
		ANTENNAMAXAREACAR 1.770800 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.148500 LAYER M2 ;
		ANTENNAMAXAREACAR 11.182300 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.066300 LAYER M3 ;
		ANTENNAMAXAREACAR 13.994800 LAYER M3 ;
	END DM[9]

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 2.575 18.890 2.725 ;
			LAYER M3 ;
			RECT 18.710 2.575 18.890 2.725 ;
			LAYER M1 ;
			RECT 18.710 2.575 18.890 2.725 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[0]

	PIN D[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 25.775 18.890 25.925 ;
			LAYER M3 ;
			RECT 18.710 25.775 18.890 25.925 ;
			LAYER M2 ;
			RECT 18.710 25.775 18.890 25.925 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[10]

	PIN D[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 28.095 18.890 28.245 ;
			LAYER M3 ;
			RECT 18.710 28.095 18.890 28.245 ;
			LAYER M2 ;
			RECT 18.710 28.095 18.890 28.245 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[11]

	PIN D[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 30.415 18.890 30.565 ;
			LAYER M1 ;
			RECT 18.710 30.415 18.890 30.565 ;
			LAYER M2 ;
			RECT 18.710 30.415 18.890 30.565 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[12]

	PIN D[13]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 32.735 18.890 32.885 ;
			LAYER M2 ;
			RECT 18.710 32.735 18.890 32.885 ;
			LAYER M1 ;
			RECT 18.710 32.735 18.890 32.885 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[13]

	PIN D[14]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 35.055 18.890 35.205 ;
			LAYER M3 ;
			RECT 18.710 35.055 18.890 35.205 ;
			LAYER M1 ;
			RECT 18.710 35.055 18.890 35.205 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[14]

	PIN D[15]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 37.375 18.890 37.525 ;
			LAYER M3 ;
			RECT 18.710 37.375 18.890 37.525 ;
			LAYER M1 ;
			RECT 18.710 37.375 18.890 37.525 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[15]

	PIN D[16]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 39.695 18.890 39.845 ;
			LAYER M1 ;
			RECT 18.710 39.695 18.890 39.845 ;
			LAYER M2 ;
			RECT 18.710 39.695 18.890 39.845 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[16]

	PIN D[17]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 42.015 18.890 42.165 ;
			LAYER M2 ;
			RECT 18.710 42.015 18.890 42.165 ;
			LAYER M1 ;
			RECT 18.710 42.015 18.890 42.165 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[17]

	PIN D[18]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 44.335 18.890 44.485 ;
			LAYER M3 ;
			RECT 18.710 44.335 18.890 44.485 ;
			LAYER M2 ;
			RECT 18.710 44.335 18.890 44.485 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[18]

	PIN D[19]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 46.655 18.890 46.805 ;
			LAYER M1 ;
			RECT 18.710 46.655 18.890 46.805 ;
			LAYER M3 ;
			RECT 18.710 46.655 18.890 46.805 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[19]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 4.895 18.890 5.045 ;
			LAYER M2 ;
			RECT 18.710 4.895 18.890 5.045 ;
			LAYER M1 ;
			RECT 18.710 4.895 18.890 5.045 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[1]

	PIN D[20]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 48.975 18.890 49.125 ;
			LAYER M1 ;
			RECT 18.710 48.975 18.890 49.125 ;
			LAYER M2 ;
			RECT 18.710 48.975 18.890 49.125 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[20]

	PIN D[21]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 51.295 18.890 51.445 ;
			LAYER M1 ;
			RECT 18.710 51.295 18.890 51.445 ;
			LAYER M2 ;
			RECT 18.710 51.295 18.890 51.445 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[21]

	PIN D[22]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 53.615 18.890 53.765 ;
			LAYER M1 ;
			RECT 18.710 53.615 18.890 53.765 ;
			LAYER M2 ;
			RECT 18.710 53.615 18.890 53.765 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[22]

	PIN D[23]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 55.935 18.890 56.085 ;
			LAYER M3 ;
			RECT 18.710 55.935 18.890 56.085 ;
			LAYER M1 ;
			RECT 18.710 55.935 18.890 56.085 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[23]

	PIN D[24]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 58.255 18.890 58.405 ;
			LAYER M1 ;
			RECT 18.710 58.255 18.890 58.405 ;
			LAYER M3 ;
			RECT 18.710 58.255 18.890 58.405 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[24]

	PIN D[25]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 80.575 18.890 80.725 ;
			LAYER M3 ;
			RECT 18.710 80.575 18.890 80.725 ;
			LAYER M2 ;
			RECT 18.710 80.575 18.890 80.725 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[25]

	PIN D[26]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 82.895 18.890 83.045 ;
			LAYER M3 ;
			RECT 18.710 82.895 18.890 83.045 ;
			LAYER M1 ;
			RECT 18.710 82.895 18.890 83.045 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[26]

	PIN D[27]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 85.215 18.890 85.365 ;
			LAYER M1 ;
			RECT 18.710 85.215 18.890 85.365 ;
			LAYER M3 ;
			RECT 18.710 85.215 18.890 85.365 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[27]

	PIN D[28]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 87.535 18.890 87.685 ;
			LAYER M1 ;
			RECT 18.710 87.535 18.890 87.685 ;
			LAYER M3 ;
			RECT 18.710 87.535 18.890 87.685 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[28]

	PIN D[29]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 89.855 18.890 90.005 ;
			LAYER M3 ;
			RECT 18.710 89.855 18.890 90.005 ;
			LAYER M1 ;
			RECT 18.710 89.855 18.890 90.005 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[29]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 7.215 18.890 7.365 ;
			LAYER M2 ;
			RECT 18.710 7.215 18.890 7.365 ;
			LAYER M3 ;
			RECT 18.710 7.215 18.890 7.365 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[2]

	PIN D[30]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 92.175 18.890 92.325 ;
			LAYER M1 ;
			RECT 18.710 92.175 18.890 92.325 ;
			LAYER M2 ;
			RECT 18.710 92.175 18.890 92.325 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[30]

	PIN D[31]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 94.495 18.890 94.645 ;
			LAYER M1 ;
			RECT 18.710 94.495 18.890 94.645 ;
			LAYER M2 ;
			RECT 18.710 94.495 18.890 94.645 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[31]

	PIN D[32]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 96.815 18.890 96.965 ;
			LAYER M3 ;
			RECT 18.710 96.815 18.890 96.965 ;
			LAYER M2 ;
			RECT 18.710 96.815 18.890 96.965 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[32]

	PIN D[33]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 99.135 18.890 99.285 ;
			LAYER M1 ;
			RECT 18.710 99.135 18.890 99.285 ;
			LAYER M3 ;
			RECT 18.710 99.135 18.890 99.285 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[33]

	PIN D[34]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 101.455 18.890 101.605 ;
			LAYER M1 ;
			RECT 18.710 101.455 18.890 101.605 ;
			LAYER M2 ;
			RECT 18.710 101.455 18.890 101.605 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[34]

	PIN D[35]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 103.775 18.890 103.925 ;
			LAYER M1 ;
			RECT 18.710 103.775 18.890 103.925 ;
			LAYER M3 ;
			RECT 18.710 103.775 18.890 103.925 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[35]

	PIN D[36]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 106.095 18.890 106.245 ;
			LAYER M2 ;
			RECT 18.710 106.095 18.890 106.245 ;
			LAYER M3 ;
			RECT 18.710 106.095 18.890 106.245 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[36]

	PIN D[37]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 108.415 18.890 108.565 ;
			LAYER M2 ;
			RECT 18.710 108.415 18.890 108.565 ;
			LAYER M1 ;
			RECT 18.710 108.415 18.890 108.565 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[37]

	PIN D[38]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 110.735 18.890 110.885 ;
			LAYER M1 ;
			RECT 18.710 110.735 18.890 110.885 ;
			LAYER M3 ;
			RECT 18.710 110.735 18.890 110.885 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[38]

	PIN D[39]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 113.055 18.890 113.205 ;
			LAYER M2 ;
			RECT 18.710 113.055 18.890 113.205 ;
			LAYER M1 ;
			RECT 18.710 113.055 18.890 113.205 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[39]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 9.535 18.890 9.685 ;
			LAYER M2 ;
			RECT 18.710 9.535 18.890 9.685 ;
			LAYER M1 ;
			RECT 18.710 9.535 18.890 9.685 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[3]

	PIN D[40]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 115.375 18.890 115.525 ;
			LAYER M1 ;
			RECT 18.710 115.375 18.890 115.525 ;
			LAYER M3 ;
			RECT 18.710 115.375 18.890 115.525 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[40]

	PIN D[41]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 117.695 18.890 117.845 ;
			LAYER M2 ;
			RECT 18.710 117.695 18.890 117.845 ;
			LAYER M3 ;
			RECT 18.710 117.695 18.890 117.845 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[41]

	PIN D[42]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 120.015 18.890 120.165 ;
			LAYER M1 ;
			RECT 18.710 120.015 18.890 120.165 ;
			LAYER M2 ;
			RECT 18.710 120.015 18.890 120.165 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[42]

	PIN D[43]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 122.335 18.890 122.485 ;
			LAYER M2 ;
			RECT 18.710 122.335 18.890 122.485 ;
			LAYER M1 ;
			RECT 18.710 122.335 18.890 122.485 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[43]

	PIN D[44]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 124.655 18.890 124.805 ;
			LAYER M1 ;
			RECT 18.710 124.655 18.890 124.805 ;
			LAYER M3 ;
			RECT 18.710 124.655 18.890 124.805 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[44]

	PIN D[45]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 126.975 18.890 127.125 ;
			LAYER M3 ;
			RECT 18.710 126.975 18.890 127.125 ;
			LAYER M1 ;
			RECT 18.710 126.975 18.890 127.125 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[45]

	PIN D[46]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 129.295 18.890 129.445 ;
			LAYER M3 ;
			RECT 18.710 129.295 18.890 129.445 ;
			LAYER M1 ;
			RECT 18.710 129.295 18.890 129.445 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[46]

	PIN D[47]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 131.615 18.890 131.765 ;
			LAYER M3 ;
			RECT 18.710 131.615 18.890 131.765 ;
			LAYER M2 ;
			RECT 18.710 131.615 18.890 131.765 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[47]

	PIN D[48]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 133.935 18.890 134.085 ;
			LAYER M1 ;
			RECT 18.710 133.935 18.890 134.085 ;
			LAYER M2 ;
			RECT 18.710 133.935 18.890 134.085 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[48]

	PIN D[49]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 136.255 18.890 136.405 ;
			LAYER M3 ;
			RECT 18.710 136.255 18.890 136.405 ;
			LAYER M2 ;
			RECT 18.710 136.255 18.890 136.405 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[49]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 11.855 18.890 12.005 ;
			LAYER M3 ;
			RECT 18.710 11.855 18.890 12.005 ;
			LAYER M1 ;
			RECT 18.710 11.855 18.890 12.005 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 14.175 18.890 14.325 ;
			LAYER M2 ;
			RECT 18.710 14.175 18.890 14.325 ;
			LAYER M1 ;
			RECT 18.710 14.175 18.890 14.325 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 16.495 18.890 16.645 ;
			LAYER M3 ;
			RECT 18.710 16.495 18.890 16.645 ;
			LAYER M1 ;
			RECT 18.710 16.495 18.890 16.645 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 18.815 18.890 18.965 ;
			LAYER M3 ;
			RECT 18.710 18.815 18.890 18.965 ;
			LAYER M2 ;
			RECT 18.710 18.815 18.890 18.965 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[7]

	PIN D[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 21.135 18.890 21.285 ;
			LAYER M2 ;
			RECT 18.710 21.135 18.890 21.285 ;
			LAYER M1 ;
			RECT 18.710 21.135 18.890 21.285 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[8]

	PIN D[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 23.455 18.890 23.605 ;
			LAYER M2 ;
			RECT 18.710 23.455 18.890 23.605 ;
			LAYER M3 ;
			RECT 18.710 23.455 18.890 23.605 ;
		END
		ANTENNAGATEAREA 0.009600 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.128000 LAYER M1 ;
		ANTENNAMAXAREACAR 13.335900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.677100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009600 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.119700 LAYER M2 ;
		ANTENNAMAXAREACAR 16.148400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.354200 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009600 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.085300 LAYER M3 ;
		ANTENNAMAXAREACAR 21.638000 LAYER M3 ;
	END D[9]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 1.930 18.890 2.080 ;
			LAYER M2 ;
			RECT 18.710 1.930 18.890 2.080 ;
			LAYER M3 ;
			RECT 18.710 1.930 18.890 2.080 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[0]

	PIN Q[10]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 25.130 18.890 25.280 ;
			LAYER M1 ;
			RECT 18.710 25.130 18.890 25.280 ;
			LAYER M3 ;
			RECT 18.710 25.130 18.890 25.280 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[10]

	PIN Q[11]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 27.450 18.890 27.600 ;
			LAYER M3 ;
			RECT 18.710 27.450 18.890 27.600 ;
			LAYER M1 ;
			RECT 18.710 27.450 18.890 27.600 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[11]

	PIN Q[12]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 29.770 18.890 29.920 ;
			LAYER M1 ;
			RECT 18.710 29.770 18.890 29.920 ;
			LAYER M2 ;
			RECT 18.710 29.770 18.890 29.920 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[12]

	PIN Q[13]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 32.090 18.890 32.240 ;
			LAYER M2 ;
			RECT 18.710 32.090 18.890 32.240 ;
			LAYER M1 ;
			RECT 18.710 32.090 18.890 32.240 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[13]

	PIN Q[14]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 34.410 18.890 34.560 ;
			LAYER M1 ;
			RECT 18.710 34.410 18.890 34.560 ;
			LAYER M3 ;
			RECT 18.710 34.410 18.890 34.560 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[14]

	PIN Q[15]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 36.730 18.890 36.880 ;
			LAYER M1 ;
			RECT 18.710 36.730 18.890 36.880 ;
			LAYER M3 ;
			RECT 18.710 36.730 18.890 36.880 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[15]

	PIN Q[16]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 39.050 18.890 39.200 ;
			LAYER M3 ;
			RECT 18.710 39.050 18.890 39.200 ;
			LAYER M2 ;
			RECT 18.710 39.050 18.890 39.200 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[16]

	PIN Q[17]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 41.370 18.890 41.520 ;
			LAYER M2 ;
			RECT 18.710 41.370 18.890 41.520 ;
			LAYER M3 ;
			RECT 18.710 41.370 18.890 41.520 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[17]

	PIN Q[18]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 43.690 18.890 43.840 ;
			LAYER M1 ;
			RECT 18.710 43.690 18.890 43.840 ;
			LAYER M3 ;
			RECT 18.710 43.690 18.890 43.840 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[18]

	PIN Q[19]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 46.010 18.890 46.160 ;
			LAYER M3 ;
			RECT 18.710 46.010 18.890 46.160 ;
			LAYER M1 ;
			RECT 18.710 46.010 18.890 46.160 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[19]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 4.250 18.890 4.400 ;
			LAYER M2 ;
			RECT 18.710 4.250 18.890 4.400 ;
			LAYER M3 ;
			RECT 18.710 4.250 18.890 4.400 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[1]

	PIN Q[20]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 48.330 18.890 48.480 ;
			LAYER M2 ;
			RECT 18.710 48.330 18.890 48.480 ;
			LAYER M3 ;
			RECT 18.710 48.330 18.890 48.480 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[20]

	PIN Q[21]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 50.650 18.890 50.800 ;
			LAYER M3 ;
			RECT 18.710 50.650 18.890 50.800 ;
			LAYER M1 ;
			RECT 18.710 50.650 18.890 50.800 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[21]

	PIN Q[22]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 52.970 18.890 53.120 ;
			LAYER M2 ;
			RECT 18.710 52.970 18.890 53.120 ;
			LAYER M3 ;
			RECT 18.710 52.970 18.890 53.120 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[22]

	PIN Q[23]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 55.290 18.890 55.440 ;
			LAYER M1 ;
			RECT 18.710 55.290 18.890 55.440 ;
			LAYER M2 ;
			RECT 18.710 55.290 18.890 55.440 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[23]

	PIN Q[24]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 57.610 18.890 57.760 ;
			LAYER M2 ;
			RECT 18.710 57.610 18.890 57.760 ;
			LAYER M1 ;
			RECT 18.710 57.610 18.890 57.760 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[24]

	PIN Q[25]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 79.930 18.890 80.080 ;
			LAYER M1 ;
			RECT 18.710 79.930 18.890 80.080 ;
			LAYER M3 ;
			RECT 18.710 79.930 18.890 80.080 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[25]

	PIN Q[26]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 82.250 18.890 82.400 ;
			LAYER M3 ;
			RECT 18.710 82.250 18.890 82.400 ;
			LAYER M1 ;
			RECT 18.710 82.250 18.890 82.400 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[26]

	PIN Q[27]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 84.570 18.890 84.720 ;
			LAYER M2 ;
			RECT 18.710 84.570 18.890 84.720 ;
			LAYER M1 ;
			RECT 18.710 84.570 18.890 84.720 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[27]

	PIN Q[28]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 86.890 18.890 87.040 ;
			LAYER M2 ;
			RECT 18.710 86.890 18.890 87.040 ;
			LAYER M1 ;
			RECT 18.710 86.890 18.890 87.040 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[28]

	PIN Q[29]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 89.210 18.890 89.360 ;
			LAYER M2 ;
			RECT 18.710 89.210 18.890 89.360 ;
			LAYER M3 ;
			RECT 18.710 89.210 18.890 89.360 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[29]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 6.570 18.890 6.720 ;
			LAYER M2 ;
			RECT 18.710 6.570 18.890 6.720 ;
			LAYER M1 ;
			RECT 18.710 6.570 18.890 6.720 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[2]

	PIN Q[30]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 91.530 18.890 91.680 ;
			LAYER M1 ;
			RECT 18.710 91.530 18.890 91.680 ;
			LAYER M2 ;
			RECT 18.710 91.530 18.890 91.680 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[30]

	PIN Q[31]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 93.850 18.890 94.000 ;
			LAYER M2 ;
			RECT 18.710 93.850 18.890 94.000 ;
			LAYER M1 ;
			RECT 18.710 93.850 18.890 94.000 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[31]

	PIN Q[32]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 96.170 18.890 96.320 ;
			LAYER M3 ;
			RECT 18.710 96.170 18.890 96.320 ;
			LAYER M2 ;
			RECT 18.710 96.170 18.890 96.320 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[32]

	PIN Q[33]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 98.490 18.890 98.640 ;
			LAYER M2 ;
			RECT 18.710 98.490 18.890 98.640 ;
			LAYER M3 ;
			RECT 18.710 98.490 18.890 98.640 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[33]

	PIN Q[34]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 100.810 18.890 100.960 ;
			LAYER M2 ;
			RECT 18.710 100.810 18.890 100.960 ;
			LAYER M1 ;
			RECT 18.710 100.810 18.890 100.960 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[34]

	PIN Q[35]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 103.130 18.890 103.280 ;
			LAYER M3 ;
			RECT 18.710 103.130 18.890 103.280 ;
			LAYER M1 ;
			RECT 18.710 103.130 18.890 103.280 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[35]

	PIN Q[36]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 105.450 18.890 105.600 ;
			LAYER M3 ;
			RECT 18.710 105.450 18.890 105.600 ;
			LAYER M1 ;
			RECT 18.710 105.450 18.890 105.600 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[36]

	PIN Q[37]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 107.770 18.890 107.920 ;
			LAYER M2 ;
			RECT 18.710 107.770 18.890 107.920 ;
			LAYER M1 ;
			RECT 18.710 107.770 18.890 107.920 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[37]

	PIN Q[38]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 110.090 18.890 110.240 ;
			LAYER M3 ;
			RECT 18.710 110.090 18.890 110.240 ;
			LAYER M2 ;
			RECT 18.710 110.090 18.890 110.240 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[38]

	PIN Q[39]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 112.410 18.890 112.560 ;
			LAYER M1 ;
			RECT 18.710 112.410 18.890 112.560 ;
			LAYER M3 ;
			RECT 18.710 112.410 18.890 112.560 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[39]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 8.890 18.890 9.040 ;
			LAYER M1 ;
			RECT 18.710 8.890 18.890 9.040 ;
			LAYER M2 ;
			RECT 18.710 8.890 18.890 9.040 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[3]

	PIN Q[40]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 114.730 18.890 114.880 ;
			LAYER M2 ;
			RECT 18.710 114.730 18.890 114.880 ;
			LAYER M3 ;
			RECT 18.710 114.730 18.890 114.880 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[40]

	PIN Q[41]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 117.050 18.890 117.200 ;
			LAYER M3 ;
			RECT 18.710 117.050 18.890 117.200 ;
			LAYER M1 ;
			RECT 18.710 117.050 18.890 117.200 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[41]

	PIN Q[42]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 119.370 18.890 119.520 ;
			LAYER M1 ;
			RECT 18.710 119.370 18.890 119.520 ;
			LAYER M2 ;
			RECT 18.710 119.370 18.890 119.520 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[42]

	PIN Q[43]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 121.690 18.890 121.840 ;
			LAYER M2 ;
			RECT 18.710 121.690 18.890 121.840 ;
			LAYER M3 ;
			RECT 18.710 121.690 18.890 121.840 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[43]

	PIN Q[44]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 124.010 18.890 124.160 ;
			LAYER M2 ;
			RECT 18.710 124.010 18.890 124.160 ;
			LAYER M1 ;
			RECT 18.710 124.010 18.890 124.160 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[44]

	PIN Q[45]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 126.330 18.890 126.480 ;
			LAYER M3 ;
			RECT 18.710 126.330 18.890 126.480 ;
			LAYER M1 ;
			RECT 18.710 126.330 18.890 126.480 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[45]

	PIN Q[46]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 128.650 18.890 128.800 ;
			LAYER M2 ;
			RECT 18.710 128.650 18.890 128.800 ;
			LAYER M3 ;
			RECT 18.710 128.650 18.890 128.800 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[46]

	PIN Q[47]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 130.970 18.890 131.120 ;
			LAYER M1 ;
			RECT 18.710 130.970 18.890 131.120 ;
			LAYER M3 ;
			RECT 18.710 130.970 18.890 131.120 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[47]

	PIN Q[48]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 133.290 18.890 133.440 ;
			LAYER M2 ;
			RECT 18.710 133.290 18.890 133.440 ;
			LAYER M3 ;
			RECT 18.710 133.290 18.890 133.440 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[48]

	PIN Q[49]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 135.610 18.890 135.760 ;
			LAYER M1 ;
			RECT 18.710 135.610 18.890 135.760 ;
			LAYER M2 ;
			RECT 18.710 135.610 18.890 135.760 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[49]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 11.210 18.890 11.360 ;
			LAYER M3 ;
			RECT 18.710 11.210 18.890 11.360 ;
			LAYER M2 ;
			RECT 18.710 11.210 18.890 11.360 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 13.530 18.890 13.680 ;
			LAYER M2 ;
			RECT 18.710 13.530 18.890 13.680 ;
			LAYER M3 ;
			RECT 18.710 13.530 18.890 13.680 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 15.850 18.890 16.000 ;
			LAYER M3 ;
			RECT 18.710 15.850 18.890 16.000 ;
			LAYER M2 ;
			RECT 18.710 15.850 18.890 16.000 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 18.170 18.890 18.320 ;
			LAYER M3 ;
			RECT 18.710 18.170 18.890 18.320 ;
			LAYER M2 ;
			RECT 18.710 18.170 18.890 18.320 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[7]

	PIN Q[8]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 20.490 18.890 20.640 ;
			LAYER M1 ;
			RECT 18.710 20.490 18.890 20.640 ;
			LAYER M2 ;
			RECT 18.710 20.490 18.890 20.640 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[8]

	PIN Q[9]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 22.810 18.890 22.960 ;
			LAYER M1 ;
			RECT 18.710 22.810 18.890 22.960 ;
			LAYER M2 ;
			RECT 18.710 22.810 18.890 22.960 ;
		END
		ANTENNADIFFAREA 0.107000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.251700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNADIFFAREA 0.107000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.226000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA2 ;
		ANTENNADIFFAREA 0.107000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.093500 LAYER M3 ;
	END Q[9]

	PIN RTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 77.605 18.890 77.755 ;
			LAYER M3 ;
			RECT 18.710 77.605 18.890 77.755 ;
			LAYER M1 ;
			RECT 18.710 77.605 18.890 77.755 ;
		END
		ANTENNAGATEAREA 0.009000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.068500 LAYER M1 ;
		ANTENNAMAXAREACAR 3.266700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.722200 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.183700 LAYER M2 ;
		ANTENNAMAXAREACAR 129.367000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.444400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.126300 LAYER M3 ;
		ANTENNAMAXAREACAR 132.367000 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 2.166700 LAYER VIA3 ;
		ANTENNAGATEAREA 0.009000 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 7.277400 LAYER M4 ;
		ANTENNAMAXAREACAR 821.700000 LAYER M4 ;
	END RTSEL[0]

	PIN RTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 77.935 18.890 78.085 ;
			LAYER M2 ;
			RECT 18.710 77.935 18.890 78.085 ;
			LAYER M1 ;
			RECT 18.710 77.935 18.890 78.085 ;
		END
		ANTENNAGATEAREA 0.009000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.068500 LAYER M1 ;
		ANTENNAMAXAREACAR 3.266700 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.722200 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 1.183700 LAYER M2 ;
		ANTENNAMAXAREACAR 129.367000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.032500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.444400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.126300 LAYER M3 ;
		ANTENNAMAXAREACAR 132.367000 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 2.166700 LAYER VIA3 ;
		ANTENNAGATEAREA 0.009000 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 7.277400 LAYER M4 ;
		ANTENNAMAXAREACAR 821.700000 LAYER M4 ;
	END RTSEL[1]

	PIN SD
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 73.735 18.890 73.885 ;
			LAYER M1 ;
			RECT 18.710 73.735 18.890 73.885 ;
			LAYER M3 ;
			RECT 18.710 73.735 18.890 73.885 ;
		END
		ANTENNAGATEAREA 0.037800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.204300 LAYER M1 ;
		ANTENNAMAXAREACAR 1.638900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.172000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.037800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.229800 LAYER M2 ;
		ANTENNAMAXAREACAR 2.938100 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.037800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.541400 LAYER M3 ;
		ANTENNAMAXAREACAR 14.542300 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 0.515900 LAYER VIA3 ;
		ANTENNAGATEAREA 0.037800 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 7.283800 LAYER M4 ;
		ANTENNAMAXAREACAR 142.553000 LAYER M4 ;
	END SD

	PIN SLP
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 18.710 73.345 18.890 73.495 ;
			LAYER M2 ;
			RECT 18.710 73.345 18.890 73.495 ;
			LAYER M3 ;
			RECT 18.710 73.345 18.890 73.495 ;
		END
		ANTENNAGATEAREA 0.037800 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.171600 LAYER M1 ;
		ANTENNAMAXAREACAR 0.688900 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.172000 LAYER VIA1 ;
		ANTENNAGATEAREA 0.037800 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.209700 LAYER M2 ;
		ANTENNAMAXAREACAR 2.153400 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.026000 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.343900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.037800 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.321200 LAYER M3 ;
		ANTENNAMAXAREACAR 4.765900 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 0.515900 LAYER VIA3 ;
		ANTENNAGATEAREA 0.037800 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 12.153600 LAYER M4 ;
		ANTENNAMAXAREACAR 197.254000 LAYER M4 ;
	END SLP

	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M4 ;
			RECT 0.000 2.815 18.505 3.105 ;
			LAYER M4 ;
			RECT 0.000 5.135 18.505 5.425 ;
			LAYER M4 ;
			RECT 0.000 7.455 18.505 7.745 ;
			LAYER M4 ;
			RECT 0.000 9.775 18.505 10.065 ;
			LAYER M4 ;
			RECT 0.000 12.095 18.505 12.385 ;
			LAYER M4 ;
			RECT 0.000 14.415 18.505 14.705 ;
			LAYER M4 ;
			RECT 0.000 16.735 18.505 17.025 ;
			LAYER M4 ;
			RECT 0.000 19.055 18.505 19.345 ;
			LAYER M4 ;
			RECT 0.000 21.375 18.505 21.665 ;
			LAYER M4 ;
			RECT 0.000 23.695 18.505 23.985 ;
			LAYER M4 ;
			RECT 0.000 26.015 18.505 26.305 ;
			LAYER M4 ;
			RECT 0.000 28.335 18.505 28.625 ;
			LAYER M4 ;
			RECT 0.000 30.655 18.505 30.945 ;
			LAYER M4 ;
			RECT 0.000 32.975 18.505 33.265 ;
			LAYER M4 ;
			RECT 0.000 35.295 18.505 35.585 ;
			LAYER M4 ;
			RECT 0.000 37.615 18.505 37.905 ;
			LAYER M4 ;
			RECT 0.000 39.935 18.505 40.225 ;
			LAYER M4 ;
			RECT 0.000 42.255 18.505 42.545 ;
			LAYER M4 ;
			RECT 0.000 44.575 18.505 44.865 ;
			LAYER M4 ;
			RECT 0.000 46.895 18.505 47.185 ;
			LAYER M4 ;
			RECT 0.000 49.215 18.505 49.505 ;
			LAYER M4 ;
			RECT 0.000 51.535 18.505 51.825 ;
			LAYER M4 ;
			RECT 0.000 53.855 18.505 54.145 ;
			LAYER M4 ;
			RECT 0.000 56.175 18.505 56.465 ;
			LAYER M4 ;
			RECT 0.000 58.495 18.505 58.785 ;
			LAYER M4 ;
			RECT 0.000 62.135 18.555 62.555 ;
			LAYER M4 ;
			RECT 0.000 65.405 18.555 65.825 ;
			LAYER M4 ;
			RECT 0.000 72.805 18.555 73.225 ;
			LAYER M4 ;
			RECT 0.000 76.330 18.555 76.750 ;
			LAYER M4 ;
			RECT 0.000 80.815 18.505 81.105 ;
			LAYER M4 ;
			RECT 0.000 83.135 18.505 83.425 ;
			LAYER M4 ;
			RECT 0.000 85.455 18.505 85.745 ;
			LAYER M4 ;
			RECT 0.000 87.775 18.505 88.065 ;
			LAYER M4 ;
			RECT 0.000 90.095 18.505 90.385 ;
			LAYER M4 ;
			RECT 0.000 92.415 18.505 92.705 ;
			LAYER M4 ;
			RECT 0.000 94.735 18.505 95.025 ;
			LAYER M4 ;
			RECT 0.000 97.055 18.505 97.345 ;
			LAYER M4 ;
			RECT 0.000 99.375 18.505 99.665 ;
			LAYER M4 ;
			RECT 0.000 101.695 18.505 101.985 ;
			LAYER M4 ;
			RECT 0.000 104.015 18.505 104.305 ;
			LAYER M4 ;
			RECT 0.000 106.335 18.505 106.625 ;
			LAYER M4 ;
			RECT 0.000 108.655 18.505 108.945 ;
			LAYER M4 ;
			RECT 0.000 110.975 18.505 111.265 ;
			LAYER M4 ;
			RECT 0.000 113.295 18.505 113.585 ;
			LAYER M4 ;
			RECT 0.000 115.615 18.505 115.905 ;
			LAYER M4 ;
			RECT 0.000 117.935 18.505 118.225 ;
			LAYER M4 ;
			RECT 0.000 120.255 18.505 120.545 ;
			LAYER M4 ;
			RECT 0.000 122.575 18.505 122.865 ;
			LAYER M4 ;
			RECT 0.000 124.895 18.505 125.185 ;
			LAYER M4 ;
			RECT 0.000 127.215 18.505 127.505 ;
			LAYER M4 ;
			RECT 0.000 129.535 18.505 129.825 ;
			LAYER M4 ;
			RECT 0.000 131.855 18.505 132.145 ;
			LAYER M4 ;
			RECT 0.000 134.175 18.505 134.465 ;
			LAYER M4 ;
			RECT 0.000 136.495 18.505 136.785 ;
		END
	END VDD

	PIN VSS
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M4 ;
			RECT 0.000 0.885 18.505 1.175 ;
			LAYER M4 ;
			RECT 0.000 3.205 18.505 3.495 ;
			LAYER M4 ;
			RECT 0.000 5.525 18.505 5.815 ;
			LAYER M4 ;
			RECT 0.000 7.845 18.505 8.135 ;
			LAYER M4 ;
			RECT 0.000 10.165 18.505 10.455 ;
			LAYER M4 ;
			RECT 0.000 12.485 18.505 12.775 ;
			LAYER M4 ;
			RECT 0.000 14.805 18.505 15.095 ;
			LAYER M4 ;
			RECT 0.000 17.125 18.505 17.415 ;
			LAYER M4 ;
			RECT 0.000 19.445 18.505 19.735 ;
			LAYER M4 ;
			RECT 0.000 21.765 18.505 22.055 ;
			LAYER M4 ;
			RECT 0.000 24.085 18.505 24.375 ;
			LAYER M4 ;
			RECT 0.000 26.405 18.505 26.695 ;
			LAYER M4 ;
			RECT 0.000 28.725 18.505 29.015 ;
			LAYER M4 ;
			RECT 0.000 31.045 18.505 31.335 ;
			LAYER M4 ;
			RECT 0.000 33.365 18.505 33.655 ;
			LAYER M4 ;
			RECT 0.000 35.685 18.505 35.975 ;
			LAYER M4 ;
			RECT 0.000 38.005 18.505 38.295 ;
			LAYER M4 ;
			RECT 0.000 40.325 18.505 40.615 ;
			LAYER M4 ;
			RECT 0.000 42.645 18.505 42.935 ;
			LAYER M4 ;
			RECT 0.000 44.965 18.505 45.255 ;
			LAYER M4 ;
			RECT 0.000 47.285 18.505 47.575 ;
			LAYER M4 ;
			RECT 0.000 49.605 18.505 49.895 ;
			LAYER M4 ;
			RECT 0.000 51.925 18.505 52.215 ;
			LAYER M4 ;
			RECT 0.000 54.245 18.505 54.535 ;
			LAYER M4 ;
			RECT 0.000 56.565 18.505 56.855 ;
			LAYER M4 ;
			RECT 0.000 63.715 18.555 64.135 ;
			LAYER M4 ;
			RECT 0.000 67.830 18.555 68.250 ;
			LAYER M4 ;
			RECT 0.000 70.785 18.555 71.205 ;
			LAYER M4 ;
			RECT 0.000 74.175 18.555 74.595 ;
			LAYER M4 ;
			RECT 0.000 78.885 18.505 79.175 ;
			LAYER M4 ;
			RECT 0.000 81.205 18.505 81.495 ;
			LAYER M4 ;
			RECT 0.000 83.525 18.505 83.815 ;
			LAYER M4 ;
			RECT 0.000 85.845 18.505 86.135 ;
			LAYER M4 ;
			RECT 0.000 88.165 18.505 88.455 ;
			LAYER M4 ;
			RECT 0.000 90.485 18.505 90.775 ;
			LAYER M4 ;
			RECT 0.000 92.805 18.505 93.095 ;
			LAYER M4 ;
			RECT 0.000 95.125 18.505 95.415 ;
			LAYER M4 ;
			RECT 0.000 97.445 18.505 97.735 ;
			LAYER M4 ;
			RECT 0.000 99.765 18.505 100.055 ;
			LAYER M4 ;
			RECT 0.000 102.085 18.505 102.375 ;
			LAYER M4 ;
			RECT 0.000 104.405 18.505 104.695 ;
			LAYER M4 ;
			RECT 0.000 106.725 18.505 107.015 ;
			LAYER M4 ;
			RECT 0.000 109.045 18.505 109.335 ;
			LAYER M4 ;
			RECT 0.000 111.365 18.505 111.655 ;
			LAYER M4 ;
			RECT 0.000 113.685 18.505 113.975 ;
			LAYER M4 ;
			RECT 0.000 116.005 18.505 116.295 ;
			LAYER M4 ;
			RECT 0.000 118.325 18.505 118.615 ;
			LAYER M4 ;
			RECT 0.000 120.645 18.505 120.935 ;
			LAYER M4 ;
			RECT 0.000 122.965 18.505 123.255 ;
			LAYER M4 ;
			RECT 0.000 125.285 18.505 125.575 ;
			LAYER M4 ;
			RECT 0.000 127.605 18.505 127.895 ;
			LAYER M4 ;
			RECT 0.000 129.925 18.505 130.215 ;
			LAYER M4 ;
			RECT 0.000 132.245 18.505 132.535 ;
			LAYER M4 ;
			RECT 0.000 134.565 18.505 134.855 ;
		END
	END VSS

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 65.440 18.890 65.590 ;
			LAYER M2 ;
			RECT 18.710 65.440 18.890 65.590 ;
			LAYER M1 ;
			RECT 18.710 65.440 18.890 65.590 ;
		END
		ANTENNAGATEAREA 0.030000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.084700 LAYER M1 ;
		ANTENNAMAXAREACAR 2.040000 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.393900 LAYER VIA1 ;
		ANTENNAGATEAREA 0.030000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.131800 LAYER M2 ;
		ANTENNAMAXAREACAR 5.010600 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.590900 LAYER VIA2 ;
		ANTENNAGATEAREA 0.030000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.828800 LAYER M3 ;
	END WEB

	PIN WEBM
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 65.900 18.890 66.050 ;
			LAYER M1 ;
			RECT 18.710 65.900 18.890 66.050 ;
			LAYER M3 ;
			RECT 18.710 65.900 18.890 66.050 ;
		END
		ANTENNAGATEAREA 0.033000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.152900 LAYER M1 ;
		ANTENNAMAXAREACAR 3.005600 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.361100 LAYER VIA1 ;
		ANTENNAGATEAREA 0.033000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.092700 LAYER M2 ;
		ANTENNAMAXAREACAR 5.066700 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.006500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 0.505600 LAYER VIA2 ;
		ANTENNAGATEAREA 0.033000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.027000 LAYER M3 ;
		ANTENNAMAXAREACAR 5.772700 LAYER M3 ;
	END WEBM

	PIN WTSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 18.710 76.850 18.890 77.000 ;
			LAYER M1 ;
			RECT 18.710 76.850 18.890 77.000 ;
			LAYER M3 ;
			RECT 18.710 76.850 18.890 77.000 ;
		END
		ANTENNAGATEAREA 0.009000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.088500 LAYER M1 ;
		ANTENNAMAXAREACAR 5.483300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.722200 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.960700 LAYER M2 ;
		ANTENNAMAXAREACAR 110.600000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.444400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.180500 LAYER M3 ;
		ANTENNAMAXAREACAR 113.600000 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 2.166700 LAYER VIA3 ;
		ANTENNAGATEAREA 0.009000 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 7.088100 LAYER M4 ;
		ANTENNAMAXAREACAR 799.264000 LAYER M4 ;
	END WTSEL[0]

	PIN WTSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 18.710 78.265 18.890 78.415 ;
			LAYER M2 ;
			RECT 18.710 78.265 18.890 78.415 ;
			LAYER M1 ;
			RECT 18.710 78.265 18.890 78.415 ;
		END
		ANTENNAGATEAREA 0.009000 LAYER M1 ;
		ANTENNADIFFAREA 0.020000 LAYER M1 ;
		ANTENNAPARTIALMETALAREA 0.088500 LAYER M1 ;
		ANTENNAMAXAREACAR 5.483300 LAYER M1 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA1 ;
		ANTENNAMAXAREACAR 0.722200 LAYER VIA1 ;
		ANTENNAGATEAREA 0.009000 LAYER M2 ;
		ANTENNADIFFAREA 0.020000 LAYER M2 ;
		ANTENNAPARTIALMETALAREA 0.960700 LAYER M2 ;
		ANTENNAMAXAREACAR 110.600000 LAYER M2 ;
		ANTENNAPARTIALCUTAREA 0.019500 LAYER VIA2 ;
		ANTENNAMAXAREACAR 1.444400 LAYER VIA2 ;
		ANTENNAGATEAREA 0.009000 LAYER M3 ;
		ANTENNADIFFAREA 0.020000 LAYER M3 ;
		ANTENNAPARTIALMETALAREA 0.180500 LAYER M3 ;
		ANTENNAMAXAREACAR 113.600000 LAYER M3 ;
		ANTENNAPARTIALCUTAREA 0.013000 LAYER VIA3 ;
		ANTENNAMAXAREACAR 2.166700 LAYER VIA3 ;
		ANTENNAGATEAREA 0.009000 LAYER M4 ;
		ANTENNADIFFAREA 0.020000 LAYER M4 ;
		ANTENNAPARTIALMETALAREA 7.088100 LAYER M4 ;
		ANTENNAMAXAREACAR 799.264000 LAYER M4 ;
	END WTSEL[1]

	OBS
		# Promoted blockages
		LAYER M1 ;
		RECT 18.710 136.795 18.890 137.670 ;
		LAYER M3 ;
		RECT 18.710 134.845 18.890 134.865 ;
		LAYER VIA3 ;
		RECT 18.710 134.845 18.890 134.865 ;
		LAYER M3 ;
		RECT 18.710 134.495 18.890 134.535 ;
		LAYER VIA3 ;
		RECT 18.710 136.815 18.890 137.670 ;
		LAYER M1 ;
		RECT 18.710 134.145 18.890 134.205 ;
		LAYER VIA3 ;
		RECT 18.710 134.495 18.890 134.535 ;
		LAYER M1 ;
		RECT 18.710 134.475 18.890 134.555 ;
		LAYER M1 ;
		RECT 18.710 121.235 18.890 121.630 ;
		LAYER VIA3 ;
		RECT 18.710 121.255 18.890 121.610 ;
		LAYER VIA3 ;
		RECT 18.710 132.525 18.890 132.545 ;
		LAYER M1 ;
		RECT 18.710 128.860 18.890 129.235 ;
		LAYER VIA3 ;
		RECT 18.710 127.885 18.890 127.905 ;
		LAYER M3 ;
		RECT 18.710 127.535 18.890 127.575 ;
		LAYER VIA3 ;
		RECT 18.710 127.535 18.890 127.575 ;
		LAYER M1 ;
		RECT 18.710 127.515 18.890 127.595 ;
		LAYER M3 ;
		RECT 18.710 127.885 18.890 127.905 ;
		LAYER M2 ;
		RECT 18.710 127.885 18.890 127.905 ;
		LAYER M2 ;
		RECT 18.710 127.205 18.890 127.225 ;
		LAYER VIA3 ;
		RECT 18.710 126.560 18.890 126.895 ;
		LAYER M3 ;
		RECT 18.710 126.560 18.890 126.895 ;
		LAYER VIA3 ;
		RECT 18.710 125.565 18.890 125.585 ;
		LAYER VIA3 ;
		RECT 18.710 122.565 18.890 122.585 ;
		LAYER VIA3 ;
		RECT 18.710 122.895 18.890 122.935 ;
		LAYER M3 ;
		RECT 18.710 122.895 18.890 122.935 ;
		LAYER M3 ;
		RECT 18.710 121.255 18.890 121.610 ;
		LAYER M2 ;
		RECT 18.710 121.255 18.890 121.610 ;
		LAYER M2 ;
		RECT 18.710 123.575 18.890 123.930 ;
		LAYER M3 ;
		RECT 18.710 123.245 18.890 123.265 ;
		LAYER M2 ;
		RECT 18.710 125.565 18.890 125.585 ;
		LAYER VIA3 ;
		RECT 18.710 125.215 18.890 125.255 ;
		LAYER M2 ;
		RECT 18.710 125.215 18.890 125.255 ;
		LAYER M3 ;
		RECT 18.710 124.885 18.890 124.905 ;
		LAYER M1 ;
		RECT 18.710 95.715 18.890 96.110 ;
		LAYER M2 ;
		RECT 18.710 100.045 18.890 100.065 ;
		LAYER M1 ;
		RECT 18.710 99.675 18.890 99.755 ;
		LAYER M2 ;
		RECT 18.710 99.365 18.890 99.385 ;
		LAYER M3 ;
		RECT 18.710 99.695 18.890 99.735 ;
		LAYER VIA3 ;
		RECT 18.710 99.695 18.890 99.735 ;
		LAYER M2 ;
		RECT 18.710 99.695 18.890 99.735 ;
		LAYER M1 ;
		RECT 18.710 108.625 18.890 108.685 ;
		LAYER M1 ;
		RECT 18.710 100.025 18.890 100.085 ;
		LAYER M1 ;
		RECT 18.710 103.340 18.890 103.715 ;
		LAYER M2 ;
		RECT 18.710 100.375 18.890 100.730 ;
		LAYER M2 ;
		RECT 18.710 89.440 18.890 89.775 ;
		LAYER M1 ;
		RECT 18.710 89.420 18.890 89.795 ;
		LAYER VIA3 ;
		RECT 18.710 90.085 18.890 90.105 ;
		LAYER M2 ;
		RECT 18.710 90.085 18.890 90.105 ;
		LAYER M3 ;
		RECT 18.710 98.055 18.890 98.410 ;
		LAYER M3 ;
		RECT 18.710 97.725 18.890 97.745 ;
		LAYER M1 ;
		RECT 18.710 97.355 18.890 97.435 ;
		LAYER M1 ;
		RECT 18.710 98.700 18.890 99.075 ;
		LAYER M1 ;
		RECT 18.710 98.035 18.890 98.430 ;
		LAYER M3 ;
		RECT 18.710 90.085 18.890 90.105 ;
		LAYER M3 ;
		RECT 18.710 98.720 18.890 99.055 ;
		LAYER M1 ;
		RECT 18.710 90.395 18.890 90.475 ;
		LAYER M3 ;
		RECT 18.710 89.440 18.890 89.775 ;
		LAYER VIA3 ;
		RECT 18.710 89.440 18.890 89.775 ;
		LAYER M1 ;
		RECT 18.710 90.065 18.890 90.125 ;
		LAYER M2 ;
		RECT 18.710 90.415 18.890 90.455 ;
		LAYER M1 ;
		RECT 18.710 90.745 18.890 90.805 ;
		LAYER M1 ;
		RECT 18.710 91.075 18.890 91.470 ;
		LAYER M3 ;
		RECT 18.710 91.760 18.890 92.095 ;
		LAYER M2 ;
		RECT 18.710 91.760 18.890 92.095 ;
		LAYER M2 ;
		RECT 18.710 92.405 18.890 92.425 ;
		LAYER M3 ;
		RECT 18.710 92.405 18.890 92.425 ;
		LAYER M1 ;
		RECT 18.710 92.385 18.890 92.445 ;
		LAYER M1 ;
		RECT 18.710 92.715 18.890 92.795 ;
		LAYER VIA3 ;
		RECT 18.710 92.735 18.890 92.775 ;
		LAYER VIA3 ;
		RECT 18.710 92.405 18.890 92.425 ;
		LAYER M2 ;
		RECT 18.710 92.735 18.890 92.775 ;
		LAYER M3 ;
		RECT 18.710 92.735 18.890 92.775 ;
		LAYER M3 ;
		RECT 18.710 93.415 18.890 93.770 ;
		LAYER M1 ;
		RECT 18.710 93.065 18.890 93.125 ;
		LAYER M1 ;
		RECT 18.710 95.035 18.890 95.115 ;
		LAYER M3 ;
		RECT 18.710 94.725 18.890 94.745 ;
		LAYER M1 ;
		RECT 18.710 93.395 18.890 93.790 ;
		LAYER M3 ;
		RECT 18.710 94.080 18.890 94.415 ;
		LAYER VIA3 ;
		RECT 18.710 94.080 18.890 94.415 ;
		LAYER M3 ;
		RECT 18.710 95.055 18.890 95.095 ;
		LAYER M3 ;
		RECT 18.710 90.415 18.890 90.455 ;
		LAYER VIA3 ;
		RECT 18.710 90.415 18.890 90.455 ;
		LAYER M1 ;
		RECT 18.710 91.740 18.890 92.115 ;
		LAYER M2 ;
		RECT 18.710 93.085 18.890 93.105 ;
		LAYER VIA3 ;
		RECT 18.710 93.085 18.890 93.105 ;
		LAYER M3 ;
		RECT 18.710 93.085 18.890 93.105 ;
		LAYER M2 ;
		RECT 18.710 93.415 18.890 93.770 ;
		LAYER VIA3 ;
		RECT 18.710 90.765 18.890 90.785 ;
		LAYER M2 ;
		RECT 18.710 90.765 18.890 90.785 ;
		LAYER M2 ;
		RECT 18.710 91.095 18.890 91.450 ;
		LAYER VIA3 ;
		RECT 18.710 91.095 18.890 91.450 ;
		LAYER M3 ;
		RECT 18.710 91.095 18.890 91.450 ;
		LAYER M3 ;
		RECT 18.710 90.765 18.890 90.785 ;
		LAYER VIA3 ;
		RECT 18.710 97.375 18.890 97.415 ;
		LAYER M2 ;
		RECT 18.710 97.045 18.890 97.065 ;
		LAYER M3 ;
		RECT 18.710 97.045 18.890 97.065 ;
		LAYER VIA3 ;
		RECT 18.710 97.045 18.890 97.065 ;
		LAYER M2 ;
		RECT 18.710 95.405 18.890 95.425 ;
		LAYER M1 ;
		RECT 18.710 95.385 18.890 95.445 ;
		LAYER VIA3 ;
		RECT 18.710 95.735 18.890 96.090 ;
		LAYER VIA3 ;
		RECT 18.710 95.405 18.890 95.425 ;
		LAYER M3 ;
		RECT 18.710 97.375 18.890 97.415 ;
		LAYER M2 ;
		RECT 18.710 95.735 18.890 96.090 ;
		LAYER M3 ;
		RECT 18.710 95.735 18.890 96.090 ;
		LAYER VIA3 ;
		RECT 18.710 96.400 18.890 96.735 ;
		LAYER M3 ;
		RECT 18.710 96.400 18.890 96.735 ;
		LAYER M2 ;
		RECT 18.710 88.775 18.890 89.130 ;
		LAYER M1 ;
		RECT 18.710 88.075 18.890 88.155 ;
		LAYER M3 ;
		RECT 18.710 88.095 18.890 88.135 ;
		LAYER VIA3 ;
		RECT 18.710 88.775 18.890 89.130 ;
		LAYER M3 ;
		RECT 18.710 85.445 18.890 85.465 ;
		LAYER M3 ;
		RECT 18.710 84.135 18.890 84.490 ;
		LAYER VIA3 ;
		RECT 18.710 84.135 18.890 84.490 ;
		LAYER M2 ;
		RECT 18.710 83.805 18.890 83.825 ;
		LAYER M2 ;
		RECT 18.710 84.135 18.890 84.490 ;
		LAYER M3 ;
		RECT 18.710 87.765 18.890 87.785 ;
		LAYER M1 ;
		RECT 18.710 87.100 18.890 87.475 ;
		LAYER M2 ;
		RECT 18.710 86.125 18.890 86.145 ;
		LAYER M1 ;
		RECT 18.710 85.755 18.890 85.835 ;
		LAYER VIA3 ;
		RECT 18.710 87.765 18.890 87.785 ;
		LAYER VIA3 ;
		RECT 18.710 87.120 18.890 87.455 ;
		LAYER M2 ;
		RECT 18.710 88.445 18.890 88.465 ;
		LAYER M3 ;
		RECT 18.710 88.445 18.890 88.465 ;
		LAYER VIA3 ;
		RECT 18.710 88.445 18.890 88.465 ;
		LAYER M2 ;
		RECT 18.710 88.095 18.890 88.135 ;
		LAYER M2 ;
		RECT 18.710 83.125 18.890 83.145 ;
		LAYER M1 ;
		RECT 18.710 83.105 18.890 83.165 ;
		LAYER M2 ;
		RECT 18.710 82.480 18.890 82.815 ;
		LAYER M3 ;
		RECT 18.710 82.480 18.890 82.815 ;
		LAYER M3 ;
		RECT 18.710 83.125 18.890 83.145 ;
		LAYER VIA3 ;
		RECT 18.710 83.125 18.890 83.145 ;
		LAYER M3 ;
		RECT 18.710 81.485 18.890 81.505 ;
		LAYER M2 ;
		RECT 18.710 81.815 18.890 82.170 ;
		LAYER M3 ;
		RECT 18.710 81.815 18.890 82.170 ;
		LAYER M2 ;
		RECT 18.710 81.485 18.890 81.505 ;
		LAYER VIA3 ;
		RECT 18.710 81.485 18.890 81.505 ;
		LAYER M1 ;
		RECT 18.710 81.465 18.890 81.525 ;
		LAYER M3 ;
		RECT 18.710 80.805 18.890 80.825 ;
		LAYER M3 ;
		RECT 18.710 79.495 18.890 79.850 ;
		LAYER VIA3 ;
		RECT 18.710 80.160 18.890 80.495 ;
		LAYER M1 ;
		RECT 18.710 80.140 18.890 80.515 ;
		LAYER M2 ;
		RECT 18.710 79.495 18.890 79.850 ;
		LAYER VIA3 ;
		RECT 18.710 81.135 18.890 81.175 ;
		LAYER M2 ;
		RECT 18.710 81.135 18.890 81.175 ;
		LAYER M1 ;
		RECT 18.710 81.115 18.890 81.195 ;
		LAYER M2 ;
		RECT 18.710 80.805 18.890 80.825 ;
		LAYER VIA3 ;
		RECT 18.710 80.805 18.890 80.825 ;
		LAYER M3 ;
		RECT 18.710 14.405 18.890 14.425 ;
		LAYER VIA3 ;
		RECT 18.710 14.405 18.890 14.425 ;
		LAYER VIA3 ;
		RECT 18.710 15.085 18.890 15.105 ;
		LAYER M1 ;
		RECT 18.710 18.380 18.890 18.755 ;
		LAYER M1 ;
		RECT 18.710 21.675 18.890 21.755 ;
		LAYER M3 ;
		RECT 18.710 22.045 18.890 22.065 ;
		LAYER VIA3 ;
		RECT 18.710 23.040 18.890 23.375 ;
		LAYER M1 ;
		RECT 18.710 42.555 18.890 42.635 ;
		LAYER VIA3 ;
		RECT 18.710 49.535 18.890 49.575 ;
		LAYER M3 ;
		RECT 18.710 49.535 18.890 49.575 ;
		LAYER VIA3 ;
		RECT 18.710 43.920 18.890 44.255 ;
		LAYER M1 ;
		RECT 18.710 44.545 18.890 44.605 ;
		LAYER VIA3 ;
		RECT 18.710 46.240 18.890 46.575 ;
		LAYER M1 ;
		RECT 18.710 47.875 18.890 48.270 ;
		LAYER M3 ;
		RECT 18.710 45.575 18.890 45.930 ;
		LAYER M1 ;
		RECT 18.710 14.715 18.890 14.795 ;
		LAYER M2 ;
		RECT 18.710 15.085 18.890 15.105 ;
		LAYER M3 ;
		RECT 18.710 15.085 18.890 15.105 ;
		LAYER VIA3 ;
		RECT 18.710 17.055 18.890 17.095 ;
		LAYER M2 ;
		RECT 18.710 16.080 18.890 16.415 ;
		LAYER M2 ;
		RECT 18.710 14.735 18.890 14.775 ;
		LAYER M1 ;
		RECT 18.710 17.035 18.890 17.115 ;
		LAYER M3 ;
		RECT 18.710 17.405 18.890 17.425 ;
		LAYER M1 ;
		RECT 18.710 17.385 18.890 17.445 ;
		LAYER M2 ;
		RECT 18.710 19.375 18.890 19.415 ;
		LAYER M3 ;
		RECT 18.710 19.045 18.890 19.065 ;
		LAYER VIA3 ;
		RECT 18.710 18.400 18.890 18.735 ;
		LAYER M3 ;
		RECT 18.710 18.400 18.890 18.735 ;
		LAYER VIA3 ;
		RECT 18.710 19.045 18.890 19.065 ;
		LAYER VIA3 ;
		RECT 18.710 19.375 18.890 19.415 ;
		LAYER M2 ;
		RECT 18.710 20.720 18.890 21.055 ;
		LAYER VIA3 ;
		RECT 18.710 20.720 18.890 21.055 ;
		LAYER M3 ;
		RECT 18.710 21.365 18.890 21.385 ;
		LAYER M3 ;
		RECT 18.710 19.375 18.890 19.415 ;
		LAYER M3 ;
		RECT 18.710 19.725 18.890 19.745 ;
		LAYER VIA3 ;
		RECT 18.710 19.725 18.890 19.745 ;
		LAYER M2 ;
		RECT 18.710 23.685 18.890 23.705 ;
		LAYER M3 ;
		RECT 18.710 24.695 18.890 25.050 ;
		LAYER VIA3 ;
		RECT 18.710 24.695 18.890 25.050 ;
		LAYER M3 ;
		RECT 18.710 28.325 18.890 28.345 ;
		LAYER M1 ;
		RECT 18.710 35.265 18.890 35.325 ;
		LAYER M3 ;
		RECT 18.710 33.975 18.890 34.330 ;
		LAYER VIA3 ;
		RECT 18.710 32.965 18.890 32.985 ;
		LAYER M1 ;
		RECT 18.710 36.275 18.890 36.670 ;
		LAYER VIA3 ;
		RECT 18.710 36.295 18.890 36.650 ;
		LAYER VIA3 ;
		RECT 18.710 35.285 18.890 35.305 ;
		LAYER VIA3 ;
		RECT 18.710 39.925 18.890 39.945 ;
		LAYER M2 ;
		RECT 18.710 39.925 18.890 39.945 ;
		LAYER VIA3 ;
		RECT 18.710 40.255 18.890 40.295 ;
		LAYER M1 ;
		RECT 18.710 38.595 18.890 38.990 ;
		LAYER VIA3 ;
		RECT 18.710 40.605 18.890 40.625 ;
		LAYER M1 ;
		RECT 18.710 40.915 18.890 41.310 ;
		LAYER VIA3 ;
		RECT 18.710 41.600 18.890 41.935 ;
		LAYER M3 ;
		RECT 18.710 42.575 18.890 42.615 ;
		LAYER M3 ;
		RECT 18.710 36.960 18.890 37.295 ;
		LAYER VIA3 ;
		RECT 18.710 36.960 18.890 37.295 ;
		LAYER VIA3 ;
		RECT 18.710 29.005 18.890 29.025 ;
		LAYER M3 ;
		RECT 18.710 16.725 18.890 16.745 ;
		LAYER M1 ;
		RECT 18.710 16.705 18.890 16.765 ;
		LAYER M2 ;
		RECT 18.710 17.055 18.890 17.095 ;
		LAYER M3 ;
		RECT 18.710 16.080 18.890 16.415 ;
		LAYER M3 ;
		RECT 18.710 17.055 18.890 17.095 ;
		LAYER M2 ;
		RECT 18.710 17.735 18.890 18.090 ;
		LAYER M3 ;
		RECT 18.710 17.735 18.890 18.090 ;
		LAYER VIA3 ;
		RECT 18.710 17.735 18.890 18.090 ;
		LAYER M2 ;
		RECT 18.710 17.405 18.890 17.425 ;
		LAYER M1 ;
		RECT 18.710 17.715 18.890 18.110 ;
		LAYER VIA3 ;
		RECT 18.710 17.405 18.890 17.425 ;
		LAYER M1 ;
		RECT 18.710 19.355 18.890 19.435 ;
		LAYER M2 ;
		RECT 18.710 19.045 18.890 19.065 ;
		LAYER M1 ;
		RECT 18.710 19.025 18.890 19.085 ;
		LAYER M2 ;
		RECT 18.710 18.400 18.890 18.735 ;
		LAYER M2 ;
		RECT 18.710 16.725 18.890 16.745 ;
		LAYER VIA3 ;
		RECT 18.710 16.725 18.890 16.745 ;
		LAYER M1 ;
		RECT 18.710 16.060 18.890 16.435 ;
		LAYER VIA3 ;
		RECT 18.710 16.080 18.890 16.415 ;
		LAYER M1 ;
		RECT 18.710 88.425 18.890 88.485 ;
		LAYER M2 ;
		RECT 18.710 87.120 18.890 87.455 ;
		LAYER M3 ;
		RECT 18.710 87.120 18.890 87.455 ;
		LAYER M1 ;
		RECT 18.710 86.435 18.890 86.830 ;
		LAYER M1 ;
		RECT 18.710 88.755 18.890 89.150 ;
		LAYER M3 ;
		RECT 18.710 80.160 18.890 80.495 ;
		LAYER M3 ;
		RECT 18.710 81.135 18.890 81.175 ;
		LAYER M3 ;
		RECT 18.710 83.455 18.890 83.495 ;
		LAYER M1 ;
		RECT 18.710 83.435 18.890 83.515 ;
		LAYER M1 ;
		RECT 18.710 79.475 18.890 79.870 ;
		LAYER M3 ;
		RECT 18.710 79.165 18.890 79.185 ;
		LAYER M2 ;
		RECT 18.710 79.165 18.890 79.185 ;
		LAYER M3 ;
		RECT 18.710 78.495 18.890 78.855 ;
		LAYER VIA3 ;
		RECT 18.710 79.495 18.890 79.850 ;
		LAYER VIA3 ;
		RECT 18.710 78.495 18.890 78.855 ;
		LAYER M2 ;
		RECT 18.710 78.495 18.890 78.855 ;
		LAYER M3 ;
		RECT 18.710 88.775 18.890 89.130 ;
		LAYER M1 ;
		RECT 18.710 78.475 18.890 78.875 ;
		LAYER M1 ;
		RECT 18.710 78.145 18.890 78.205 ;
		LAYER M3 ;
		RECT 18.710 77.835 18.890 77.855 ;
		LAYER M3 ;
		RECT 18.710 78.165 18.890 78.185 ;
		LAYER VIA3 ;
		RECT 18.710 78.165 18.890 78.185 ;
		LAYER M2 ;
		RECT 18.710 78.165 18.890 78.185 ;
		LAYER M3 ;
		RECT 18.710 74.295 18.890 75.990 ;
		LAYER M2 ;
		RECT 18.710 74.295 18.890 75.990 ;
		LAYER VIA3 ;
		RECT 18.710 72.440 18.890 72.590 ;
		LAYER M2 ;
		RECT 18.710 71.010 18.890 71.030 ;
		LAYER M3 ;
		RECT 18.710 70.550 18.890 70.700 ;
		LAYER M1 ;
		RECT 18.710 66.110 18.890 69.160 ;
		LAYER VIA3 ;
		RECT 18.710 66.130 18.890 69.140 ;
		LAYER M3 ;
		RECT 18.710 65.670 18.890 65.820 ;
		LAYER M3 ;
		RECT 18.710 62.330 18.890 65.360 ;
		LAYER VIA3 ;
		RECT 18.710 65.670 18.890 65.820 ;
		LAYER M1 ;
		RECT 18.710 65.650 18.890 65.840 ;
		LAYER M2 ;
		RECT 18.710 96.400 18.890 96.735 ;
		LAYER M1 ;
		RECT 18.710 97.025 18.890 97.085 ;
		LAYER M1 ;
		RECT 18.710 99.345 18.890 99.405 ;
		LAYER M2 ;
		RECT 18.710 101.040 18.890 101.375 ;
		LAYER M2 ;
		RECT 18.710 95.055 18.890 95.095 ;
		LAYER M3 ;
		RECT 18.710 110.320 18.890 110.655 ;
		LAYER VIA3 ;
		RECT 18.710 110.320 18.890 110.655 ;
		LAYER M1 ;
		RECT 18.710 57.820 18.890 58.195 ;
		LAYER M3 ;
		RECT 18.710 54.525 18.890 54.545 ;
		LAYER M3 ;
		RECT 18.710 54.175 18.890 54.215 ;
		LAYER M3 ;
		RECT 18.710 52.535 18.890 52.890 ;
		LAYER M3 ;
		RECT 18.710 58.485 18.890 58.505 ;
		LAYER VIA3 ;
		RECT 18.710 52.205 18.890 52.225 ;
		LAYER M2 ;
		RECT 18.710 52.535 18.890 52.890 ;
		LAYER M1 ;
		RECT 18.710 52.185 18.890 52.245 ;
		LAYER M2 ;
		RECT 18.710 14.405 18.890 14.425 ;
		LAYER M3 ;
		RECT 18.710 13.760 18.890 14.095 ;
		LAYER VIA3 ;
		RECT 18.710 13.760 18.890 14.095 ;
		LAYER VIA3 ;
		RECT 18.710 13.095 18.890 13.450 ;
		LAYER M3 ;
		RECT 18.710 10.775 18.890 11.130 ;
		LAYER VIA3 ;
		RECT 18.710 10.445 18.890 10.465 ;
		LAYER M3 ;
		RECT 18.710 10.445 18.890 10.465 ;
		LAYER M2 ;
		RECT 18.710 9.120 18.890 9.455 ;
		LAYER M3 ;
		RECT 18.710 9.120 18.890 9.455 ;
		LAYER M1 ;
		RECT 18.710 13.075 18.890 13.470 ;
		LAYER M1 ;
		RECT 18.710 10.075 18.890 10.155 ;
		LAYER M2 ;
		RECT 18.710 15.415 18.890 15.770 ;
		LAYER M2 ;
		RECT 18.710 8.455 18.890 8.810 ;
		LAYER M3 ;
		RECT 18.710 8.455 18.890 8.810 ;
		LAYER VIA3 ;
		RECT 18.710 8.455 18.890 8.810 ;
		LAYER M3 ;
		RECT 18.710 15.415 18.890 15.770 ;
		LAYER M3 ;
		RECT 18.710 7.775 18.890 7.815 ;
		LAYER VIA3 ;
		RECT 18.710 8.125 18.890 8.145 ;
		LAYER M1 ;
		RECT 18.710 8.435 18.890 8.830 ;
		LAYER M3 ;
		RECT 18.710 10.095 18.890 10.135 ;
		LAYER M2 ;
		RECT 18.710 10.095 18.890 10.135 ;
		LAYER M2 ;
		RECT 18.710 9.765 18.890 9.785 ;
		LAYER M1 ;
		RECT 18.710 9.745 18.890 9.805 ;
		LAYER M1 ;
		RECT 18.710 3.465 18.890 3.525 ;
		LAYER M1 ;
		RECT 18.710 2.140 18.890 2.515 ;
		LAYER M1 ;
		RECT 18.710 1.475 18.890 1.870 ;
		LAYER M2 ;
		RECT 18.710 0.000 18.890 0.855 ;
		LAYER M2 ;
		RECT 18.710 3.485 18.890 3.505 ;
		LAYER VIA3 ;
		RECT 18.710 1.165 18.890 1.185 ;
		LAYER M3 ;
		RECT 18.710 1.165 18.890 1.185 ;
		LAYER VIA3 ;
		RECT 18.710 3.485 18.890 3.505 ;
		LAYER VIA3 ;
		RECT 18.710 0.000 18.890 0.855 ;
		LAYER M1 ;
		RECT 18.710 0.000 18.890 0.875 ;
		LAYER M3 ;
		RECT 18.710 0.000 18.890 0.855 ;
		LAYER M1 ;
		RECT 18.710 1.145 18.890 1.205 ;
		LAYER M2 ;
		RECT 18.710 1.495 18.890 1.850 ;
		LAYER VIA3 ;
		RECT 18.710 1.495 18.890 1.850 ;
		LAYER M3 ;
		RECT 18.710 1.495 18.890 1.850 ;
		LAYER M2 ;
		RECT 18.710 1.165 18.890 1.185 ;
		LAYER M2 ;
		RECT 18.710 3.135 18.890 3.175 ;
		LAYER M2 ;
		RECT 18.710 2.805 18.890 2.825 ;
		LAYER M3 ;
		RECT 18.710 2.805 18.890 2.825 ;
		LAYER VIA3 ;
		RECT 18.710 2.805 18.890 2.825 ;
		LAYER M1 ;
		RECT 18.710 3.115 18.890 3.195 ;
		LAYER M1 ;
		RECT 18.710 5.435 18.890 5.515 ;
		LAYER VIA3 ;
		RECT 18.710 5.455 18.890 5.495 ;
		LAYER M2 ;
		RECT 18.710 5.455 18.890 5.495 ;
		LAYER M3 ;
		RECT 18.710 5.455 18.890 5.495 ;
		LAYER M2 ;
		RECT 18.710 5.125 18.890 5.145 ;
		LAYER M3 ;
		RECT 18.710 5.125 18.890 5.145 ;
		LAYER M1 ;
		RECT 18.710 6.115 18.890 6.510 ;
		LAYER VIA3 ;
		RECT 18.710 5.125 18.890 5.145 ;
		LAYER M1 ;
		RECT 18.710 5.105 18.890 5.165 ;
		LAYER M3 ;
		RECT 18.710 3.135 18.890 3.175 ;
		LAYER M3 ;
		RECT 18.710 3.485 18.890 3.505 ;
		LAYER M1 ;
		RECT 18.710 3.795 18.890 4.190 ;
		LAYER M1 ;
		RECT 18.710 2.785 18.890 2.845 ;
		LAYER M3 ;
		RECT 18.710 2.160 18.890 2.495 ;
		LAYER M2 ;
		RECT 18.710 2.160 18.890 2.495 ;
		LAYER VIA3 ;
		RECT 18.710 2.160 18.890 2.495 ;
		LAYER VIA3 ;
		RECT 18.710 3.135 18.890 3.175 ;
		LAYER M2 ;
		RECT 18.710 3.815 18.890 4.170 ;
		LAYER M3 ;
		RECT 18.710 3.815 18.890 4.170 ;
		LAYER VIA3 ;
		RECT 18.710 3.815 18.890 4.170 ;
		LAYER M2 ;
		RECT 18.710 4.480 18.890 4.815 ;
		LAYER M3 ;
		RECT 18.710 4.480 18.890 4.815 ;
		LAYER VIA3 ;
		RECT 18.710 4.480 18.890 4.815 ;
		LAYER M1 ;
		RECT 18.710 4.460 18.890 4.835 ;
		LAYER M1 ;
		RECT 18.710 135.820 18.890 136.195 ;
		LAYER M2 ;
		RECT 18.710 133.520 18.890 133.855 ;
		LAYER M2 ;
		RECT 18.710 134.165 18.890 134.185 ;
		LAYER M3 ;
		RECT 18.710 120.575 18.890 120.615 ;
		LAYER M1 ;
		RECT 18.710 120.555 18.890 120.635 ;
		LAYER M2 ;
		RECT 18.710 120.245 18.890 120.265 ;
		LAYER M1 ;
		RECT 18.710 120.225 18.890 120.285 ;
		LAYER VIA3 ;
		RECT 18.710 120.575 18.890 120.615 ;
		LAYER M2 ;
		RECT 18.710 120.575 18.890 120.615 ;
		LAYER M3 ;
		RECT 18.710 119.600 18.890 119.935 ;
		LAYER M2 ;
		RECT 18.710 119.600 18.890 119.935 ;
		LAYER VIA3 ;
		RECT 18.710 119.600 18.890 119.935 ;
		LAYER M2 ;
		RECT 18.710 107.005 18.890 107.025 ;
		LAYER M1 ;
		RECT 18.710 106.985 18.890 107.045 ;
		LAYER M2 ;
		RECT 18.710 107.335 18.890 107.690 ;
		LAYER M3 ;
		RECT 18.710 107.335 18.890 107.690 ;
		LAYER M3 ;
		RECT 18.710 107.005 18.890 107.025 ;
		LAYER VIA3 ;
		RECT 18.710 107.005 18.890 107.025 ;
		LAYER M2 ;
		RECT 18.710 108.000 18.890 108.335 ;
		LAYER M1 ;
		RECT 18.710 104.995 18.890 105.390 ;
		LAYER M2 ;
		RECT 18.710 104.685 18.890 104.705 ;
		LAYER M2 ;
		RECT 18.710 110.965 18.890 110.985 ;
		LAYER M1 ;
		RECT 18.710 110.945 18.890 111.005 ;
		LAYER M1 ;
		RECT 18.710 111.275 18.890 111.355 ;
		LAYER M3 ;
		RECT 18.710 110.965 18.890 110.985 ;
		LAYER VIA3 ;
		RECT 18.710 110.965 18.890 110.985 ;
		LAYER M1 ;
		RECT 18.710 111.955 18.890 112.350 ;
		LAYER VIA3 ;
		RECT 18.710 111.645 18.890 111.665 ;
		LAYER M1 ;
		RECT 18.710 111.625 18.890 111.685 ;
		LAYER M3 ;
		RECT 18.710 111.975 18.890 112.330 ;
		LAYER VIA3 ;
		RECT 18.710 111.975 18.890 112.330 ;
		LAYER M2 ;
		RECT 18.710 106.655 18.890 106.695 ;
		LAYER M2 ;
		RECT 18.710 105.680 18.890 106.015 ;
		LAYER M3 ;
		RECT 18.710 105.015 18.890 105.370 ;
		LAYER VIA3 ;
		RECT 18.710 105.015 18.890 105.370 ;
		LAYER M1 ;
		RECT 18.710 105.660 18.890 106.035 ;
		LAYER M3 ;
		RECT 18.710 108.975 18.890 109.015 ;
		LAYER M2 ;
		RECT 18.710 108.975 18.890 109.015 ;
		LAYER VIA3 ;
		RECT 18.710 108.975 18.890 109.015 ;
		LAYER M1 ;
		RECT 18.710 108.955 18.890 109.035 ;
		LAYER M2 ;
		RECT 18.710 109.325 18.890 109.345 ;
		LAYER M3 ;
		RECT 18.710 109.325 18.890 109.345 ;
		LAYER M2 ;
		RECT 18.710 108.645 18.890 108.665 ;
		LAYER M2 ;
		RECT 18.710 109.655 18.890 110.010 ;
		LAYER M1 ;
		RECT 18.710 109.635 18.890 110.030 ;
		LAYER M2 ;
		RECT 18.710 110.320 18.890 110.655 ;
		LAYER M1 ;
		RECT 18.710 110.300 18.890 110.675 ;
		LAYER VIA3 ;
		RECT 18.710 109.655 18.890 110.010 ;
		LAYER M3 ;
		RECT 18.710 109.655 18.890 110.010 ;
		LAYER VIA3 ;
		RECT 18.710 108.000 18.890 108.335 ;
		LAYER VIA3 ;
		RECT 18.710 106.325 18.890 106.345 ;
		LAYER M2 ;
		RECT 18.710 106.325 18.890 106.345 ;
		LAYER M3 ;
		RECT 18.710 103.360 18.890 103.695 ;
		LAYER VIA3 ;
		RECT 18.710 103.360 18.890 103.695 ;
		LAYER M2 ;
		RECT 18.710 103.360 18.890 103.695 ;
		LAYER M3 ;
		RECT 18.710 104.005 18.890 104.025 ;
		LAYER VIA3 ;
		RECT 18.710 104.005 18.890 104.025 ;
		LAYER M2 ;
		RECT 18.710 101.685 18.890 101.705 ;
		LAYER M3 ;
		RECT 18.710 104.685 18.890 104.705 ;
		LAYER M1 ;
		RECT 18.710 104.665 18.890 104.725 ;
		LAYER VIA3 ;
		RECT 18.710 104.685 18.890 104.705 ;
		LAYER M2 ;
		RECT 18.710 102.015 18.890 102.055 ;
		LAYER VIA3 ;
		RECT 18.710 101.685 18.890 101.705 ;
		LAYER M1 ;
		RECT 18.710 109.305 18.890 109.365 ;
		LAYER M2 ;
		RECT 18.710 116.285 18.890 116.305 ;
		LAYER M3 ;
		RECT 18.710 116.285 18.890 116.305 ;
		LAYER M1 ;
		RECT 18.710 115.915 18.890 115.995 ;
		LAYER VIA3 ;
		RECT 18.710 112.640 18.890 112.975 ;
		LAYER M3 ;
		RECT 18.710 112.640 18.890 112.975 ;
		LAYER VIA3 ;
		RECT 18.710 109.325 18.890 109.345 ;
		LAYER M3 ;
		RECT 18.710 118.605 18.890 118.625 ;
		LAYER VIA3 ;
		RECT 18.710 118.935 18.890 119.290 ;
		LAYER M1 ;
		RECT 18.710 113.265 18.890 113.325 ;
		LAYER M2 ;
		RECT 18.710 113.285 18.890 113.305 ;
		LAYER M1 ;
		RECT 18.710 115.585 18.890 115.645 ;
		LAYER VIA3 ;
		RECT 18.710 113.285 18.890 113.305 ;
		LAYER M2 ;
		RECT 18.710 113.615 18.890 113.655 ;
		LAYER M1 ;
		RECT 18.710 116.265 18.890 116.325 ;
		LAYER VIA3 ;
		RECT 18.710 116.285 18.890 116.305 ;
		LAYER M2 ;
		RECT 18.710 116.615 18.890 116.970 ;
		LAYER VIA3 ;
		RECT 18.710 117.280 18.890 117.615 ;
		LAYER M3 ;
		RECT 18.710 117.280 18.890 117.615 ;
		LAYER M1 ;
		RECT 18.710 114.275 18.890 114.670 ;
		LAYER M2 ;
		RECT 18.710 114.295 18.890 114.650 ;
		LAYER M3 ;
		RECT 18.710 113.965 18.890 113.985 ;
		LAYER VIA3 ;
		RECT 18.710 114.960 18.890 115.295 ;
		LAYER M3 ;
		RECT 18.710 136.815 18.890 137.670 ;
		LAYER M2 ;
		RECT 18.710 124.885 18.890 124.905 ;
		LAYER VIA3 ;
		RECT 18.710 124.240 18.890 124.575 ;
		LAYER M3 ;
		RECT 18.710 132.175 18.890 132.215 ;
		LAYER M2 ;
		RECT 18.710 132.175 18.890 132.215 ;
		LAYER M1 ;
		RECT 18.710 132.155 18.890 132.235 ;
		LAYER M3 ;
		RECT 18.710 131.845 18.890 131.865 ;
		LAYER VIA3 ;
		RECT 18.710 132.175 18.890 132.215 ;
		LAYER M1 ;
		RECT 18.710 129.505 18.890 129.565 ;
		LAYER M1 ;
		RECT 18.710 127.865 18.890 127.925 ;
		LAYER M2 ;
		RECT 18.710 126.560 18.890 126.895 ;
		LAYER M3 ;
		RECT 18.710 125.565 18.890 125.585 ;
		LAYER M2 ;
		RECT 18.710 120.925 18.890 120.945 ;
		LAYER M3 ;
		RECT 18.710 120.925 18.890 120.945 ;
		LAYER VIA3 ;
		RECT 18.710 120.925 18.890 120.945 ;
		LAYER M1 ;
		RECT 18.710 120.905 18.890 120.965 ;
		LAYER M3 ;
		RECT 18.710 121.920 18.890 122.255 ;
		LAYER M2 ;
		RECT 18.710 136.815 18.890 137.670 ;
		LAYER M2 ;
		RECT 18.710 135.175 18.890 135.530 ;
		LAYER M3 ;
		RECT 18.710 135.840 18.890 136.175 ;
		LAYER VIA3 ;
		RECT 18.710 135.175 18.890 135.530 ;
		LAYER M1 ;
		RECT 18.710 135.155 18.890 135.550 ;
		LAYER M3 ;
		RECT 18.710 135.175 18.890 135.530 ;
		LAYER M1 ;
		RECT 18.710 136.465 18.890 136.525 ;
		LAYER M2 ;
		RECT 18.710 136.485 18.890 136.505 ;
		LAYER M3 ;
		RECT 18.710 136.485 18.890 136.505 ;
		LAYER M2 ;
		RECT 18.710 135.840 18.890 136.175 ;
		LAYER VIA3 ;
		RECT 18.710 136.485 18.890 136.505 ;
		LAYER VIA3 ;
		RECT 18.710 135.840 18.890 136.175 ;
		LAYER VIA3 ;
		RECT 18.710 7.775 18.890 7.815 ;
		LAYER VIA3 ;
		RECT 18.710 133.520 18.890 133.855 ;
		LAYER M1 ;
		RECT 18.710 133.500 18.890 133.875 ;
		LAYER M2 ;
		RECT 18.710 134.845 18.890 134.865 ;
		LAYER M1 ;
		RECT 18.710 134.825 18.890 134.885 ;
		LAYER M2 ;
		RECT 18.710 134.495 18.890 134.535 ;
		LAYER M3 ;
		RECT 18.710 133.520 18.890 133.855 ;
		LAYER VIA3 ;
		RECT 18.710 134.165 18.890 134.185 ;
		LAYER M3 ;
		RECT 18.710 134.165 18.890 134.185 ;
		LAYER VIA3 ;
		RECT 18.710 99.365 18.890 99.385 ;
		LAYER VIA3 ;
		RECT 18.710 95.055 18.890 95.095 ;
		LAYER M2 ;
		RECT 18.710 94.725 18.890 94.745 ;
		LAYER VIA3 ;
		RECT 18.710 94.725 18.890 94.745 ;
		LAYER M1 ;
		RECT 18.710 48.540 18.890 48.915 ;
		LAYER M2 ;
		RECT 18.710 49.535 18.890 49.575 ;
		LAYER M2 ;
		RECT 18.710 49.885 18.890 49.905 ;
		LAYER M3 ;
		RECT 18.710 49.885 18.890 49.905 ;
		LAYER M2 ;
		RECT 18.710 48.560 18.890 48.895 ;
		LAYER M2 ;
		RECT 18.710 43.255 18.890 43.610 ;
		LAYER M3 ;
		RECT 18.710 43.255 18.890 43.610 ;
		LAYER VIA3 ;
		RECT 18.710 44.895 18.890 44.935 ;
		LAYER M2 ;
		RECT 18.710 44.895 18.890 44.935 ;
		LAYER VIA3 ;
		RECT 18.710 49.885 18.890 49.905 ;
		LAYER M2 ;
		RECT 18.710 87.765 18.890 87.785 ;
		LAYER M1 ;
		RECT 18.710 94.705 18.890 94.765 ;
		LAYER M1 ;
		RECT 18.710 94.060 18.890 94.435 ;
		LAYER M1 ;
		RECT 18.710 87.745 18.890 87.805 ;
		LAYER VIA3 ;
		RECT 18.710 91.760 18.890 92.095 ;
		LAYER VIA3 ;
		RECT 18.710 93.415 18.890 93.770 ;
		LAYER M2 ;
		RECT 18.710 94.080 18.890 94.415 ;
		LAYER VIA3 ;
		RECT 18.710 88.095 18.890 88.135 ;
		LAYER M2 ;
		RECT 18.710 12.415 18.890 12.455 ;
		LAYER VIA3 ;
		RECT 18.710 15.415 18.890 15.770 ;
		LAYER M1 ;
		RECT 18.710 15.395 18.890 15.790 ;
		LAYER M3 ;
		RECT 18.710 47.215 18.890 47.255 ;
		LAYER M2 ;
		RECT 18.710 47.215 18.890 47.255 ;
		LAYER M1 ;
		RECT 18.710 47.195 18.890 47.275 ;
		LAYER M2 ;
		RECT 18.710 46.885 18.890 46.905 ;
		LAYER VIA3 ;
		RECT 18.710 46.885 18.890 46.905 ;
		LAYER M3 ;
		RECT 18.710 46.885 18.890 46.905 ;
		LAYER M3 ;
		RECT 18.710 44.895 18.890 44.935 ;
		LAYER M1 ;
		RECT 18.710 47.545 18.890 47.605 ;
		LAYER M1 ;
		RECT 18.710 44.875 18.890 44.955 ;
		LAYER M2 ;
		RECT 18.710 12.765 18.890 12.785 ;
		LAYER M1 ;
		RECT 18.710 12.745 18.890 12.805 ;
		LAYER M2 ;
		RECT 18.710 13.095 18.890 13.450 ;
		LAYER M3 ;
		RECT 18.710 13.095 18.890 13.450 ;
		LAYER VIA3 ;
		RECT 18.710 12.765 18.890 12.785 ;
		LAYER M3 ;
		RECT 18.710 12.765 18.890 12.785 ;
		LAYER M2 ;
		RECT 18.710 13.760 18.890 14.095 ;
		LAYER M3 ;
		RECT 18.710 14.735 18.890 14.775 ;
		LAYER VIA3 ;
		RECT 18.710 14.735 18.890 14.775 ;
		LAYER M1 ;
		RECT 18.710 15.065 18.890 15.125 ;
		LAYER M1 ;
		RECT 18.710 25.340 18.890 25.715 ;
		LAYER M2 ;
		RECT 18.710 42.575 18.890 42.615 ;
		LAYER M3 ;
		RECT 18.710 29.005 18.890 29.025 ;
		LAYER M1 ;
		RECT 18.710 32.945 18.890 33.005 ;
		LAYER M1 ;
		RECT 18.710 32.300 18.890 32.675 ;
		LAYER M2 ;
		RECT 18.710 33.975 18.890 34.330 ;
		LAYER M2 ;
		RECT 18.710 43.920 18.890 44.255 ;
		LAYER M3 ;
		RECT 18.710 43.920 18.890 44.255 ;
		LAYER M1 ;
		RECT 18.710 43.900 18.890 44.275 ;
		LAYER M3 ;
		RECT 18.710 44.565 18.890 44.585 ;
		LAYER M1 ;
		RECT 18.710 45.225 18.890 45.285 ;
		LAYER M2 ;
		RECT 18.710 45.245 18.890 45.265 ;
		LAYER M3 ;
		RECT 18.710 45.245 18.890 45.265 ;
		LAYER VIA3 ;
		RECT 18.710 45.245 18.890 45.265 ;
		LAYER VIA3 ;
		RECT 18.710 45.575 18.890 45.930 ;
		LAYER M1 ;
		RECT 18.710 46.865 18.890 46.925 ;
		LAYER M1 ;
		RECT 18.710 46.220 18.890 46.595 ;
		LAYER M2 ;
		RECT 18.710 46.240 18.890 46.575 ;
		LAYER M2 ;
		RECT 18.710 45.575 18.890 45.930 ;
		LAYER M1 ;
		RECT 18.710 45.555 18.890 45.950 ;
		LAYER M1 ;
		RECT 18.710 43.235 18.890 43.630 ;
		LAYER M3 ;
		RECT 18.710 42.925 18.890 42.945 ;
		LAYER VIA3 ;
		RECT 18.710 42.925 18.890 42.945 ;
		LAYER VIA3 ;
		RECT 18.710 42.575 18.890 42.615 ;
		LAYER M2 ;
		RECT 18.710 10.445 18.890 10.465 ;
		LAYER VIA3 ;
		RECT 18.710 9.765 18.890 9.785 ;
		LAYER VIA3 ;
		RECT 18.710 9.120 18.890 9.455 ;
		LAYER M1 ;
		RECT 18.710 9.100 18.890 9.475 ;
		LAYER M3 ;
		RECT 18.710 9.765 18.890 9.785 ;
		LAYER VIA3 ;
		RECT 18.710 10.095 18.890 10.135 ;
		LAYER M2 ;
		RECT 18.710 7.775 18.890 7.815 ;
		LAYER M3 ;
		RECT 18.710 8.125 18.890 8.145 ;
		LAYER VIA3 ;
		RECT 18.710 11.440 18.890 11.775 ;
		LAYER M2 ;
		RECT 18.710 10.775 18.890 11.130 ;
		LAYER M1 ;
		RECT 18.710 7.755 18.890 7.835 ;
		LAYER M2 ;
		RECT 18.710 8.125 18.890 8.145 ;
		LAYER M2 ;
		RECT 18.710 7.445 18.890 7.465 ;
		LAYER M1 ;
		RECT 18.710 7.425 18.890 7.485 ;
		LAYER M1 ;
		RECT 18.710 6.780 18.890 7.155 ;
		LAYER M2 ;
		RECT 18.710 6.135 18.890 6.490 ;
		LAYER M3 ;
		RECT 18.710 6.800 18.890 7.135 ;
		LAYER VIA3 ;
		RECT 18.710 6.800 18.890 7.135 ;
		LAYER M1 ;
		RECT 18.710 12.395 18.890 12.475 ;
		LAYER M1 ;
		RECT 18.710 132.835 18.890 133.230 ;
		LAYER M2 ;
		RECT 18.710 132.855 18.890 133.210 ;
		LAYER M1 ;
		RECT 18.710 132.505 18.890 132.565 ;
		LAYER M3 ;
		RECT 18.710 132.525 18.890 132.545 ;
		LAYER M2 ;
		RECT 18.710 132.525 18.890 132.545 ;
		LAYER VIA3 ;
		RECT 18.710 132.855 18.890 133.210 ;
		LAYER M3 ;
		RECT 18.710 132.855 18.890 133.210 ;
		LAYER M3 ;
		RECT 18.710 50.215 18.890 50.570 ;
		LAYER M2 ;
		RECT 18.710 51.855 18.890 51.895 ;
		LAYER M3 ;
		RECT 18.710 51.855 18.890 51.895 ;
		LAYER VIA3 ;
		RECT 18.710 51.855 18.890 51.895 ;
		LAYER M1 ;
		RECT 18.710 51.835 18.890 51.915 ;
		LAYER M1 ;
		RECT 18.710 50.860 18.890 51.235 ;
		LAYER VIA3 ;
		RECT 18.710 51.525 18.890 51.545 ;
		LAYER M2 ;
		RECT 18.710 51.525 18.890 51.545 ;
		LAYER M1 ;
		RECT 18.710 51.505 18.890 51.565 ;
		LAYER M3 ;
		RECT 18.710 51.525 18.890 51.545 ;
		LAYER M2 ;
		RECT 18.710 52.205 18.890 52.225 ;
		LAYER M3 ;
		RECT 18.710 52.205 18.890 52.225 ;
		LAYER M1 ;
		RECT 18.710 52.515 18.890 52.910 ;
		LAYER M3 ;
		RECT 18.710 53.200 18.890 53.535 ;
		LAYER VIA3 ;
		RECT 18.710 53.200 18.890 53.535 ;
		LAYER VIA3 ;
		RECT 18.710 52.535 18.890 52.890 ;
		LAYER M1 ;
		RECT 18.710 53.825 18.890 53.885 ;
		LAYER M2 ;
		RECT 18.710 53.845 18.890 53.865 ;
		LAYER M2 ;
		RECT 18.710 53.200 18.890 53.535 ;
		LAYER M1 ;
		RECT 18.710 53.180 18.890 53.555 ;
		LAYER M3 ;
		RECT 18.710 53.845 18.890 53.865 ;
		LAYER VIA3 ;
		RECT 18.710 53.845 18.890 53.865 ;
		LAYER M2 ;
		RECT 18.710 77.080 18.890 77.525 ;
		LAYER M3 ;
		RECT 18.710 77.080 18.890 77.525 ;
		LAYER M2 ;
		RECT 18.710 80.160 18.890 80.495 ;
		LAYER M1 ;
		RECT 18.710 79.145 18.890 79.205 ;
		LAYER VIA3 ;
		RECT 18.710 79.165 18.890 79.185 ;
		LAYER M1 ;
		RECT 18.710 77.815 18.890 77.875 ;
		LAYER VIA3 ;
		RECT 18.710 77.835 18.890 77.855 ;
		LAYER M2 ;
		RECT 18.710 77.835 18.890 77.855 ;
		LAYER M1 ;
		RECT 18.710 77.060 18.890 77.545 ;
		LAYER VIA3 ;
		RECT 18.710 77.080 18.890 77.525 ;
		LAYER M2 ;
		RECT 18.710 76.300 18.890 76.770 ;
		LAYER M3 ;
		RECT 18.710 76.300 18.890 76.770 ;
		LAYER M3 ;
		RECT 18.710 84.800 18.890 85.135 ;
		LAYER VIA3 ;
		RECT 18.710 84.800 18.890 85.135 ;
		LAYER M1 ;
		RECT 18.710 84.780 18.890 85.155 ;
		LAYER M3 ;
		RECT 18.710 83.805 18.890 83.825 ;
		LAYER M1 ;
		RECT 18.710 84.115 18.890 84.510 ;
		LAYER M2 ;
		RECT 18.710 84.800 18.890 85.135 ;
		LAYER M3 ;
		RECT 18.710 73.965 18.890 73.985 ;
		LAYER M2 ;
		RECT 18.710 73.965 18.890 73.985 ;
		LAYER VIA3 ;
		RECT 18.710 73.965 18.890 73.985 ;
		LAYER M1 ;
		RECT 18.710 73.945 18.890 74.005 ;
		LAYER M1 ;
		RECT 18.710 76.280 18.890 76.790 ;
		LAYER VIA3 ;
		RECT 18.710 76.300 18.890 76.770 ;
		LAYER VIA3 ;
		RECT 18.710 74.295 18.890 75.990 ;
		LAYER M1 ;
		RECT 18.710 72.880 18.890 73.285 ;
		LAYER M1 ;
		RECT 18.710 74.275 18.890 76.010 ;
		LAYER M2 ;
		RECT 18.710 69.910 18.890 70.240 ;
		LAYER M3 ;
		RECT 18.710 69.910 18.890 70.240 ;
		LAYER M1 ;
		RECT 18.710 71.780 18.890 72.150 ;
		LAYER M3 ;
		RECT 18.710 72.440 18.890 72.590 ;
		LAYER M2 ;
		RECT 18.710 72.440 18.890 72.590 ;
		LAYER VIA3 ;
		RECT 18.710 70.550 18.890 70.700 ;
		LAYER M2 ;
		RECT 18.710 50.880 18.890 51.215 ;
		LAYER M3 ;
		RECT 18.710 50.880 18.890 51.215 ;
		LAYER VIA3 ;
		RECT 18.710 50.880 18.890 51.215 ;
		LAYER M3 ;
		RECT 18.710 86.125 18.890 86.145 ;
		LAYER M1 ;
		RECT 18.710 86.105 18.890 86.165 ;
		LAYER M2 ;
		RECT 18.710 86.455 18.890 86.810 ;
		LAYER M3 ;
		RECT 18.710 86.455 18.890 86.810 ;
		LAYER VIA3 ;
		RECT 18.710 86.125 18.890 86.145 ;
		LAYER VIA3 ;
		RECT 18.710 86.455 18.890 86.810 ;
		LAYER M2 ;
		RECT 18.710 50.215 18.890 50.570 ;
		LAYER VIA3 ;
		RECT 18.710 50.215 18.890 50.570 ;
		LAYER M2 ;
		RECT 18.710 54.175 18.890 54.215 ;
		LAYER M1 ;
		RECT 18.710 54.155 18.890 54.235 ;
		LAYER VIA3 ;
		RECT 18.710 54.175 18.890 54.215 ;
		LAYER M3 ;
		RECT 18.710 54.855 18.890 55.210 ;
		LAYER M1 ;
		RECT 18.710 54.835 18.890 55.230 ;
		LAYER M2 ;
		RECT 18.710 57.840 18.890 58.175 ;
		LAYER VIA3 ;
		RECT 18.710 57.840 18.890 58.175 ;
		LAYER M3 ;
		RECT 18.710 57.840 18.890 58.175 ;
		LAYER M3 ;
		RECT 18.710 85.775 18.890 85.815 ;
		LAYER M2 ;
		RECT 18.710 85.775 18.890 85.815 ;
		LAYER VIA3 ;
		RECT 18.710 85.775 18.890 85.815 ;
		LAYER M1 ;
		RECT 18.710 85.425 18.890 85.485 ;
		LAYER VIA3 ;
		RECT 18.710 85.445 18.890 85.465 ;
		LAYER M2 ;
		RECT 18.710 85.445 18.890 85.465 ;
		LAYER VIA3 ;
		RECT 18.710 83.455 18.890 83.495 ;
		LAYER VIA3 ;
		RECT 18.710 83.805 18.890 83.825 ;
		LAYER M1 ;
		RECT 18.710 83.785 18.890 83.845 ;
		LAYER M1 ;
		RECT 18.710 82.460 18.890 82.835 ;
		LAYER VIA3 ;
		RECT 18.710 82.480 18.890 82.815 ;
		LAYER M2 ;
		RECT 18.710 83.455 18.890 83.495 ;
		LAYER VIA3 ;
		RECT 18.710 81.815 18.890 82.170 ;
		LAYER M1 ;
		RECT 18.710 81.795 18.890 82.190 ;
		LAYER M1 ;
		RECT 18.710 80.785 18.890 80.845 ;
		LAYER M2 ;
		RECT 18.710 54.525 18.890 54.545 ;
		LAYER VIA3 ;
		RECT 18.710 54.525 18.890 54.545 ;
		LAYER M1 ;
		RECT 18.710 54.505 18.890 54.565 ;
		LAYER VIA3 ;
		RECT 18.710 54.855 18.890 55.210 ;
		LAYER M2 ;
		RECT 18.710 54.855 18.890 55.210 ;
		LAYER M2 ;
		RECT 18.710 56.165 18.890 56.185 ;
		LAYER M1 ;
		RECT 18.710 55.500 18.890 55.875 ;
		LAYER M1 ;
		RECT 18.710 56.145 18.890 56.205 ;
		LAYER M2 ;
		RECT 18.710 56.495 18.890 56.535 ;
		LAYER M3 ;
		RECT 18.710 56.495 18.890 56.535 ;
		LAYER VIA3 ;
		RECT 18.710 56.165 18.890 56.185 ;
		LAYER VIA3 ;
		RECT 18.710 56.495 18.890 56.535 ;
		LAYER M1 ;
		RECT 18.710 56.475 18.890 56.555 ;
		LAYER M2 ;
		RECT 18.710 56.845 18.890 56.865 ;
		LAYER M3 ;
		RECT 18.710 56.845 18.890 56.865 ;
		LAYER VIA3 ;
		RECT 18.710 56.845 18.890 56.865 ;
		LAYER M1 ;
		RECT 18.710 56.825 18.890 56.885 ;
		LAYER M1 ;
		RECT 18.710 57.155 18.890 57.550 ;
		LAYER M2 ;
		RECT 18.710 57.175 18.890 57.530 ;
		LAYER M3 ;
		RECT 18.710 57.175 18.890 57.530 ;
		LAYER VIA3 ;
		RECT 18.710 57.175 18.890 57.530 ;
		LAYER VIA3 ;
		RECT 18.710 55.520 18.890 55.855 ;
		LAYER M2 ;
		RECT 18.710 55.520 18.890 55.855 ;
		LAYER M3 ;
		RECT 18.710 55.520 18.890 55.855 ;
		LAYER M3 ;
		RECT 18.710 56.165 18.890 56.185 ;
		LAYER M1 ;
		RECT 18.710 73.555 18.890 73.675 ;
		LAYER VIA3 ;
		RECT 18.710 73.575 18.890 73.655 ;
		LAYER M2 ;
		RECT 18.710 73.575 18.890 73.655 ;
		LAYER M3 ;
		RECT 18.710 73.575 18.890 73.655 ;
		LAYER M2 ;
		RECT 18.710 72.900 18.890 73.265 ;
		LAYER VIA3 ;
		RECT 18.710 72.900 18.890 73.265 ;
		LAYER M3 ;
		RECT 18.710 72.900 18.890 73.265 ;
		LAYER M1 ;
		RECT 18.710 72.420 18.890 72.610 ;
		LAYER M1 ;
		RECT 18.710 71.320 18.890 71.510 ;
		LAYER M2 ;
		RECT 18.710 71.340 18.890 71.490 ;
		LAYER VIA3 ;
		RECT 18.710 71.340 18.890 71.490 ;
		LAYER M3 ;
		RECT 18.710 71.800 18.890 72.130 ;
		LAYER M3 ;
		RECT 18.710 71.340 18.890 71.490 ;
		LAYER M1 ;
		RECT 18.710 70.990 18.890 71.050 ;
		LAYER VIA3 ;
		RECT 18.710 71.800 18.890 72.130 ;
		LAYER M2 ;
		RECT 18.710 71.800 18.890 72.130 ;
		LAYER VIA3 ;
		RECT 18.710 71.010 18.890 71.030 ;
		LAYER VIA3 ;
		RECT 18.710 69.910 18.890 70.240 ;
		LAYER M1 ;
		RECT 18.710 69.430 18.890 69.620 ;
		LAYER M3 ;
		RECT 18.710 69.450 18.890 69.600 ;
		LAYER VIA3 ;
		RECT 18.710 69.450 18.890 69.600 ;
		LAYER M2 ;
		RECT 18.710 58.815 18.890 61.030 ;
		LAYER M1 ;
		RECT 18.710 62.310 18.890 65.380 ;
		LAYER M2 ;
		RECT 18.710 62.330 18.890 65.360 ;
		LAYER M2 ;
		RECT 18.710 65.670 18.890 65.820 ;
		LAYER M2 ;
		RECT 18.710 66.130 18.890 69.140 ;
		LAYER M3 ;
		RECT 18.710 66.130 18.890 69.140 ;
		LAYER VIA3 ;
		RECT 18.710 62.330 18.890 65.360 ;
		LAYER M1 ;
		RECT 18.710 69.890 18.890 70.260 ;
		LAYER M2 ;
		RECT 18.710 70.550 18.890 70.700 ;
		LAYER M3 ;
		RECT 18.710 71.010 18.890 71.030 ;
		LAYER M2 ;
		RECT 18.710 69.450 18.890 69.600 ;
		LAYER M1 ;
		RECT 18.710 70.530 18.890 70.720 ;
		LAYER VIA3 ;
		RECT 18.710 58.815 18.890 61.030 ;
		LAYER M1 ;
		RECT 18.710 58.795 18.890 61.050 ;
		LAYER VIA3 ;
		RECT 18.710 58.485 18.890 58.505 ;
		LAYER M1 ;
		RECT 18.710 58.465 18.890 58.525 ;
		LAYER M2 ;
		RECT 18.710 58.485 18.890 58.505 ;
		LAYER M3 ;
		RECT 18.710 58.815 18.890 61.030 ;
		LAYER M1 ;
		RECT 18.710 61.320 18.890 61.380 ;
		LAYER VIA3 ;
		RECT 18.710 61.340 18.890 61.360 ;
		LAYER M3 ;
		RECT 18.710 61.340 18.890 61.360 ;
		LAYER M2 ;
		RECT 18.710 61.340 18.890 61.360 ;
		LAYER M3 ;
		RECT 18.710 61.670 18.890 61.690 ;
		LAYER M2 ;
		RECT 18.710 61.670 18.890 61.690 ;
		LAYER VIA3 ;
		RECT 18.710 61.670 18.890 61.690 ;
		LAYER M1 ;
		RECT 18.710 61.650 18.890 61.710 ;
		LAYER M3 ;
		RECT 18.710 62.000 18.890 62.020 ;
		LAYER VIA3 ;
		RECT 18.710 62.000 18.890 62.020 ;
		LAYER M2 ;
		RECT 18.710 62.000 18.890 62.020 ;
		LAYER M1 ;
		RECT 18.710 61.980 18.890 62.040 ;
		LAYER M1 ;
		RECT 18.710 131.825 18.890 131.885 ;
		LAYER M2 ;
		RECT 18.710 131.845 18.890 131.865 ;
		LAYER VIA3 ;
		RECT 18.710 131.845 18.890 131.865 ;
		LAYER M3 ;
		RECT 18.710 131.200 18.890 131.535 ;
		LAYER M1 ;
		RECT 18.710 131.180 18.890 131.555 ;
		LAYER M2 ;
		RECT 18.710 130.535 18.890 130.890 ;
		LAYER M3 ;
		RECT 18.710 130.535 18.890 130.890 ;
		LAYER VIA3 ;
		RECT 18.710 130.535 18.890 130.890 ;
		LAYER VIA3 ;
		RECT 18.710 131.200 18.890 131.535 ;
		LAYER M2 ;
		RECT 18.710 131.200 18.890 131.535 ;
		LAYER M1 ;
		RECT 18.710 130.515 18.890 130.910 ;
		LAYER VIA3 ;
		RECT 18.710 113.965 18.890 113.985 ;
		LAYER M2 ;
		RECT 18.710 113.965 18.890 113.985 ;
		LAYER M1 ;
		RECT 18.710 113.945 18.890 114.005 ;
		LAYER M1 ;
		RECT 18.710 113.595 18.890 113.675 ;
		LAYER M2 ;
		RECT 18.710 102.365 18.890 102.385 ;
		LAYER M2 ;
		RECT 18.710 97.725 18.890 97.745 ;
		LAYER M2 ;
		RECT 18.710 98.055 18.890 98.410 ;
		LAYER VIA3 ;
		RECT 18.710 98.055 18.890 98.410 ;
		LAYER VIA3 ;
		RECT 18.710 97.725 18.890 97.745 ;
		LAYER M2 ;
		RECT 18.710 127.535 18.890 127.575 ;
		LAYER M1 ;
		RECT 18.710 127.185 18.890 127.245 ;
		LAYER M3 ;
		RECT 18.710 114.295 18.890 114.650 ;
		LAYER VIA3 ;
		RECT 18.710 114.295 18.890 114.650 ;
		LAYER M4 ;
		RECT 18.505 76.850 18.555 137.670 ;
		LAYER M1 ;
		RECT 18.710 106.635 18.890 106.715 ;
		LAYER M3 ;
		RECT 18.710 106.655 18.890 106.695 ;
		LAYER M2 ;
		RECT 18.710 112.640 18.890 112.975 ;
		LAYER M2 ;
		RECT 18.710 111.645 18.890 111.665 ;
		LAYER M3 ;
		RECT 18.710 111.645 18.890 111.665 ;
		LAYER M2 ;
		RECT 18.710 111.295 18.890 111.335 ;
		LAYER M1 ;
		RECT 18.710 101.995 18.890 102.075 ;
		LAYER M3 ;
		RECT 18.710 99.365 18.890 99.385 ;
		LAYER VIA3 ;
		RECT 18.710 100.045 18.890 100.065 ;
		LAYER M3 ;
		RECT 18.710 102.365 18.890 102.385 ;
		LAYER VIA3 ;
		RECT 18.710 98.720 18.890 99.055 ;
		LAYER M2 ;
		RECT 18.710 98.720 18.890 99.055 ;
		LAYER VIA3 ;
		RECT 18.710 129.525 18.890 129.545 ;
		LAYER VIA3 ;
		RECT 18.710 128.880 18.890 129.215 ;
		LAYER M2 ;
		RECT 18.710 128.880 18.890 129.215 ;
		LAYER M3 ;
		RECT 18.710 128.880 18.890 129.215 ;
		LAYER M2 ;
		RECT 18.710 128.215 18.890 128.570 ;
		LAYER VIA3 ;
		RECT 18.710 128.215 18.890 128.570 ;
		LAYER M3 ;
		RECT 18.710 128.215 18.890 128.570 ;
		LAYER M2 ;
		RECT 18.710 129.525 18.890 129.545 ;
		LAYER M3 ;
		RECT 18.710 129.525 18.890 129.545 ;
		LAYER M1 ;
		RECT 18.710 128.195 18.890 128.590 ;
		LAYER M1 ;
		RECT 18.710 129.835 18.890 129.915 ;
		LAYER VIA3 ;
		RECT 18.710 130.205 18.890 130.225 ;
		LAYER M2 ;
		RECT 18.710 130.205 18.890 130.225 ;
		LAYER M1 ;
		RECT 18.710 130.185 18.890 130.245 ;
		LAYER VIA3 ;
		RECT 18.710 102.365 18.890 102.385 ;
		LAYER M3 ;
		RECT 18.710 108.000 18.890 108.335 ;
		LAYER M1 ;
		RECT 18.710 107.980 18.890 108.355 ;
		LAYER VIA3 ;
		RECT 18.710 108.645 18.890 108.665 ;
		LAYER M3 ;
		RECT 18.710 108.645 18.890 108.665 ;
		LAYER M1 ;
		RECT 18.710 102.345 18.890 102.405 ;
		LAYER M2 ;
		RECT 18.710 105.015 18.890 105.370 ;
		LAYER M3 ;
		RECT 18.710 105.680 18.890 106.015 ;
		LAYER VIA3 ;
		RECT 18.710 105.680 18.890 106.015 ;
		LAYER M3 ;
		RECT 18.710 106.325 18.890 106.345 ;
		LAYER M1 ;
		RECT 18.710 106.305 18.890 106.365 ;
		LAYER VIA3 ;
		RECT 18.710 106.655 18.890 106.695 ;
		LAYER VIA3 ;
		RECT 18.710 107.335 18.890 107.690 ;
		LAYER M1 ;
		RECT 18.710 107.315 18.890 107.710 ;
		LAYER M3 ;
		RECT 18.710 101.040 18.890 101.375 ;
		LAYER M1 ;
		RECT 18.710 101.020 18.890 101.395 ;
		LAYER M3 ;
		RECT 18.710 101.685 18.890 101.705 ;
		LAYER M1 ;
		RECT 18.710 101.665 18.890 101.725 ;
		LAYER M3 ;
		RECT 18.710 102.015 18.890 102.055 ;
		LAYER VIA3 ;
		RECT 18.710 102.015 18.890 102.055 ;
		LAYER VIA3 ;
		RECT 18.710 101.040 18.890 101.375 ;
		LAYER M1 ;
		RECT 18.710 100.355 18.890 100.750 ;
		LAYER M3 ;
		RECT 18.710 100.045 18.890 100.065 ;
		LAYER M3 ;
		RECT 18.710 100.375 18.890 100.730 ;
		LAYER VIA3 ;
		RECT 18.710 100.375 18.890 100.730 ;
		LAYER VIA3 ;
		RECT 18.710 121.920 18.890 122.255 ;
		LAYER M2 ;
		RECT 18.710 118.935 18.890 119.290 ;
		LAYER M3 ;
		RECT 18.710 118.935 18.890 119.290 ;
		LAYER M2 ;
		RECT 18.710 118.255 18.890 118.295 ;
		LAYER M3 ;
		RECT 18.710 118.255 18.890 118.295 ;
		LAYER VIA3 ;
		RECT 18.710 118.255 18.890 118.295 ;
		LAYER M1 ;
		RECT 18.710 118.585 18.890 118.645 ;
		LAYER M1 ;
		RECT 18.710 122.545 18.890 122.605 ;
		LAYER M2 ;
		RECT 18.710 122.565 18.890 122.585 ;
		LAYER VIA3 ;
		RECT 18.710 116.615 18.890 116.970 ;
		LAYER M3 ;
		RECT 18.710 122.565 18.890 122.585 ;
		LAYER M1 ;
		RECT 18.710 118.235 18.890 118.315 ;
		LAYER M1 ;
		RECT 18.710 118.915 18.890 119.310 ;
		LAYER M3 ;
		RECT 18.710 115.935 18.890 115.975 ;
		LAYER M1 ;
		RECT 18.710 116.595 18.890 116.990 ;
		LAYER M2 ;
		RECT 18.710 122.895 18.890 122.935 ;
		LAYER M1 ;
		RECT 18.710 122.875 18.890 122.955 ;
		LAYER M2 ;
		RECT 18.710 115.935 18.890 115.975 ;
		LAYER M3 ;
		RECT 18.710 116.615 18.890 116.970 ;
		LAYER M1 ;
		RECT 18.710 117.905 18.890 117.965 ;
		LAYER M2 ;
		RECT 18.710 117.925 18.890 117.945 ;
		LAYER M1 ;
		RECT 18.710 117.260 18.890 117.635 ;
		LAYER M2 ;
		RECT 18.710 117.280 18.890 117.615 ;
		LAYER M3 ;
		RECT 18.710 117.925 18.890 117.945 ;
		LAYER VIA3 ;
		RECT 18.710 117.925 18.890 117.945 ;
		LAYER VIA3 ;
		RECT 18.710 115.935 18.890 115.975 ;
		LAYER M1 ;
		RECT 18.710 123.225 18.890 123.285 ;
		LAYER M2 ;
		RECT 18.710 123.245 18.890 123.265 ;
		LAYER M3 ;
		RECT 18.710 120.245 18.890 120.265 ;
		LAYER M1 ;
		RECT 18.710 119.580 18.890 119.955 ;
		LAYER VIA3 ;
		RECT 18.710 118.605 18.890 118.625 ;
		LAYER M2 ;
		RECT 18.710 118.605 18.890 118.625 ;
		LAYER VIA3 ;
		RECT 18.710 120.245 18.890 120.265 ;
		LAYER M1 ;
		RECT 18.710 123.555 18.890 123.950 ;
		LAYER M3 ;
		RECT 18.710 123.575 18.890 123.930 ;
		LAYER VIA3 ;
		RECT 18.710 123.575 18.890 123.930 ;
		LAYER M1 ;
		RECT 18.710 124.865 18.890 124.925 ;
		LAYER VIA3 ;
		RECT 18.710 124.885 18.890 124.905 ;
		LAYER M2 ;
		RECT 18.710 124.240 18.890 124.575 ;
		LAYER M3 ;
		RECT 18.710 124.240 18.890 124.575 ;
		LAYER M1 ;
		RECT 18.710 124.220 18.890 124.595 ;
		LAYER M1 ;
		RECT 18.710 126.540 18.890 126.915 ;
		LAYER M2 ;
		RECT 18.710 125.895 18.890 126.250 ;
		LAYER VIA3 ;
		RECT 18.710 125.895 18.890 126.250 ;
		LAYER M3 ;
		RECT 18.710 125.895 18.890 126.250 ;
		LAYER M1 ;
		RECT 18.710 104.315 18.890 104.395 ;
		LAYER VIA3 ;
		RECT 18.710 104.335 18.890 104.375 ;
		LAYER M3 ;
		RECT 18.710 104.335 18.890 104.375 ;
		LAYER M2 ;
		RECT 18.710 104.005 18.890 104.025 ;
		LAYER M1 ;
		RECT 18.710 103.985 18.890 104.045 ;
		LAYER M3 ;
		RECT 18.710 102.695 18.890 103.050 ;
		LAYER VIA3 ;
		RECT 18.710 102.695 18.890 103.050 ;
		LAYER M2 ;
		RECT 18.710 104.335 18.890 104.375 ;
		LAYER M1 ;
		RECT 18.710 102.675 18.890 103.070 ;
		LAYER M2 ;
		RECT 18.710 102.695 18.890 103.050 ;
		LAYER M1 ;
		RECT 18.710 114.940 18.890 115.315 ;
		LAYER M2 ;
		RECT 18.710 115.605 18.890 115.625 ;
		LAYER M3 ;
		RECT 18.710 115.605 18.890 115.625 ;
		LAYER M3 ;
		RECT 18.710 113.285 18.890 113.305 ;
		LAYER VIA3 ;
		RECT 18.710 115.605 18.890 115.625 ;
		LAYER M2 ;
		RECT 18.710 114.960 18.890 115.295 ;
		LAYER M3 ;
		RECT 18.710 114.960 18.890 115.295 ;
		LAYER M2 ;
		RECT 18.710 111.975 18.890 112.330 ;
		LAYER M1 ;
		RECT 18.710 112.620 18.890 112.995 ;
		LAYER M3 ;
		RECT 18.710 127.205 18.890 127.225 ;
		LAYER M1 ;
		RECT 18.710 125.875 18.890 126.270 ;
		LAYER M3 ;
		RECT 18.710 125.215 18.890 125.255 ;
		LAYER M1 ;
		RECT 18.710 125.545 18.890 125.605 ;
		LAYER M1 ;
		RECT 18.710 125.195 18.890 125.275 ;
		LAYER VIA3 ;
		RECT 18.710 127.205 18.890 127.225 ;
		LAYER M1 ;
		RECT 18.710 28.635 18.890 28.715 ;
		LAYER M3 ;
		RECT 18.710 28.655 18.890 28.695 ;
		LAYER VIA3 ;
		RECT 18.710 28.655 18.890 28.695 ;
		LAYER VIA3 ;
		RECT 18.710 28.325 18.890 28.345 ;
		LAYER M2 ;
		RECT 18.710 28.325 18.890 28.345 ;
		LAYER M1 ;
		RECT 18.710 33.955 18.890 34.350 ;
		LAYER VIA3 ;
		RECT 18.710 33.975 18.890 34.330 ;
		LAYER M2 ;
		RECT 18.710 32.965 18.890 32.985 ;
		LAYER M3 ;
		RECT 18.710 32.965 18.890 32.985 ;
		LAYER VIA3 ;
		RECT 18.710 27.015 18.890 27.370 ;
		LAYER M2 ;
		RECT 18.710 27.015 18.890 27.370 ;
		LAYER M3 ;
		RECT 18.710 27.015 18.890 27.370 ;
		LAYER VIA3 ;
		RECT 18.710 27.680 18.890 28.015 ;
		LAYER M1 ;
		RECT 18.710 26.995 18.890 27.390 ;
		LAYER M1 ;
		RECT 18.710 26.665 18.890 26.725 ;
		LAYER M2 ;
		RECT 18.710 26.685 18.890 26.705 ;
		LAYER M3 ;
		RECT 18.710 26.685 18.890 26.705 ;
		LAYER VIA3 ;
		RECT 18.710 26.685 18.890 26.705 ;
		LAYER M1 ;
		RECT 18.710 29.315 18.890 29.710 ;
		LAYER M1 ;
		RECT 18.710 30.625 18.890 30.685 ;
		LAYER M2 ;
		RECT 18.710 29.335 18.890 29.690 ;
		LAYER VIA3 ;
		RECT 18.710 29.335 18.890 29.690 ;
		LAYER M1 ;
		RECT 18.710 29.980 18.890 30.355 ;
		LAYER M3 ;
		RECT 18.710 29.335 18.890 29.690 ;
		LAYER M2 ;
		RECT 18.710 30.000 18.890 30.335 ;
		LAYER M3 ;
		RECT 18.710 30.000 18.890 30.335 ;
		LAYER M2 ;
		RECT 18.710 30.645 18.890 30.665 ;
		LAYER M3 ;
		RECT 18.710 30.645 18.890 30.665 ;
		LAYER VIA3 ;
		RECT 18.710 30.645 18.890 30.665 ;
		LAYER VIA3 ;
		RECT 18.710 30.000 18.890 30.335 ;
		LAYER M2 ;
		RECT 18.710 28.655 18.890 28.695 ;
		LAYER M3 ;
		RECT 18.710 32.320 18.890 32.655 ;
		LAYER VIA3 ;
		RECT 18.710 32.320 18.890 32.655 ;
		LAYER M1 ;
		RECT 18.710 28.985 18.890 29.045 ;
		LAYER M2 ;
		RECT 18.710 29.005 18.890 29.025 ;
		LAYER M2 ;
		RECT 18.710 33.645 18.890 33.665 ;
		LAYER M3 ;
		RECT 18.710 33.645 18.890 33.665 ;
		LAYER VIA3 ;
		RECT 18.710 33.645 18.890 33.665 ;
		LAYER M1 ;
		RECT 18.710 33.275 18.890 33.355 ;
		LAYER M1 ;
		RECT 18.710 30.955 18.890 31.035 ;
		LAYER M2 ;
		RECT 18.710 30.975 18.890 31.015 ;
		LAYER M3 ;
		RECT 18.710 30.975 18.890 31.015 ;
		LAYER VIA3 ;
		RECT 18.710 30.975 18.890 31.015 ;
		LAYER M2 ;
		RECT 18.710 31.655 18.890 32.010 ;
		LAYER VIA3 ;
		RECT 18.710 31.655 18.890 32.010 ;
		LAYER M3 ;
		RECT 18.710 31.325 18.890 31.345 ;
		LAYER M2 ;
		RECT 18.710 32.320 18.890 32.655 ;
		LAYER VIA3 ;
		RECT 18.710 31.325 18.890 31.345 ;
		LAYER M2 ;
		RECT 18.710 31.325 18.890 31.345 ;
		LAYER M1 ;
		RECT 18.710 28.305 18.890 28.365 ;
		LAYER M2 ;
		RECT 18.710 27.680 18.890 28.015 ;
		LAYER M3 ;
		RECT 18.710 27.680 18.890 28.015 ;
		LAYER M1 ;
		RECT 18.710 27.660 18.890 28.035 ;
		LAYER M1 ;
		RECT 18.710 33.625 18.890 33.685 ;
		LAYER M2 ;
		RECT 18.710 33.295 18.890 33.335 ;
		LAYER VIA3 ;
		RECT 18.710 33.295 18.890 33.335 ;
		LAYER M1 ;
		RECT 18.710 34.620 18.890 34.995 ;
		LAYER VIA3 ;
		RECT 18.710 34.640 18.890 34.975 ;
		LAYER M1 ;
		RECT 18.710 35.595 18.890 35.675 ;
		LAYER M1 ;
		RECT 18.710 37.915 18.890 37.995 ;
		LAYER VIA3 ;
		RECT 18.710 37.935 18.890 37.975 ;
		LAYER M3 ;
		RECT 18.710 37.605 18.890 37.625 ;
		LAYER VIA3 ;
		RECT 18.710 37.605 18.890 37.625 ;
		LAYER M3 ;
		RECT 18.710 37.935 18.890 37.975 ;
		LAYER M2 ;
		RECT 18.710 37.935 18.890 37.975 ;
		LAYER M2 ;
		RECT 18.710 36.960 18.890 37.295 ;
		LAYER M1 ;
		RECT 18.710 36.940 18.890 37.315 ;
		LAYER M2 ;
		RECT 18.710 36.295 18.890 36.650 ;
		LAYER M3 ;
		RECT 18.710 36.295 18.890 36.650 ;
		LAYER M2 ;
		RECT 18.710 35.965 18.890 35.985 ;
		LAYER M1 ;
		RECT 18.710 35.945 18.890 36.005 ;
		LAYER M2 ;
		RECT 18.710 35.615 18.890 35.655 ;
		LAYER M3 ;
		RECT 18.710 35.615 18.890 35.655 ;
		LAYER VIA3 ;
		RECT 18.710 35.965 18.890 35.985 ;
		LAYER M3 ;
		RECT 18.710 35.965 18.890 35.985 ;
		LAYER VIA3 ;
		RECT 18.710 35.615 18.890 35.655 ;
		LAYER M3 ;
		RECT 18.710 23.040 18.890 23.375 ;
		LAYER M3 ;
		RECT 18.710 20.720 18.890 21.055 ;
		LAYER M1 ;
		RECT 18.710 19.705 18.890 19.765 ;
		LAYER M1 ;
		RECT 18.710 20.700 18.890 21.075 ;
		LAYER M1 ;
		RECT 18.710 21.345 18.890 21.405 ;
		LAYER M2 ;
		RECT 18.710 21.695 18.890 21.735 ;
		LAYER VIA3 ;
		RECT 18.710 21.695 18.890 21.735 ;
		LAYER M2 ;
		RECT 18.710 21.365 18.890 21.385 ;
		LAYER M2 ;
		RECT 18.710 22.045 18.890 22.065 ;
		LAYER VIA3 ;
		RECT 18.710 21.365 18.890 21.385 ;
		LAYER M3 ;
		RECT 18.710 21.695 18.890 21.735 ;
		LAYER M1 ;
		RECT 18.710 20.035 18.890 20.430 ;
		LAYER VIA3 ;
		RECT 18.710 20.055 18.890 20.410 ;
		LAYER M2 ;
		RECT 18.710 20.055 18.890 20.410 ;
		LAYER M2 ;
		RECT 18.710 19.725 18.890 19.745 ;
		LAYER M3 ;
		RECT 18.710 20.055 18.890 20.410 ;
		LAYER VIA3 ;
		RECT 18.710 22.045 18.890 22.065 ;
		LAYER M1 ;
		RECT 18.710 22.025 18.890 22.085 ;
		LAYER VIA3 ;
		RECT 18.710 22.375 18.890 22.730 ;
		LAYER M1 ;
		RECT 18.710 22.355 18.890 22.750 ;
		LAYER M2 ;
		RECT 18.710 22.375 18.890 22.730 ;
		LAYER M3 ;
		RECT 18.710 22.375 18.890 22.730 ;
		LAYER M1 ;
		RECT 18.710 26.315 18.890 26.395 ;
		LAYER VIA3 ;
		RECT 18.710 26.335 18.890 26.375 ;
		LAYER VIA3 ;
		RECT 18.710 25.360 18.890 25.695 ;
		LAYER M1 ;
		RECT 18.710 25.985 18.890 26.045 ;
		LAYER M2 ;
		RECT 18.710 26.335 18.890 26.375 ;
		LAYER M3 ;
		RECT 18.710 26.335 18.890 26.375 ;
		LAYER M1 ;
		RECT 18.710 24.675 18.890 25.070 ;
		LAYER M2 ;
		RECT 18.710 24.695 18.890 25.050 ;
		LAYER VIA3 ;
		RECT 18.710 39.280 18.890 39.615 ;
		LAYER M3 ;
		RECT 18.710 41.600 18.890 41.935 ;
		LAYER M2 ;
		RECT 18.710 41.600 18.890 41.935 ;
		LAYER M1 ;
		RECT 18.710 41.580 18.890 41.955 ;
		LAYER M1 ;
		RECT 18.710 42.225 18.890 42.285 ;
		LAYER VIA3 ;
		RECT 18.710 42.245 18.890 42.265 ;
		LAYER M2 ;
		RECT 18.710 42.245 18.890 42.265 ;
		LAYER M3 ;
		RECT 18.710 42.245 18.890 42.265 ;
		LAYER M3 ;
		RECT 18.710 26.005 18.890 26.025 ;
		LAYER M2 ;
		RECT 18.710 26.005 18.890 26.025 ;
		LAYER M2 ;
		RECT 18.710 25.360 18.890 25.695 ;
		LAYER M3 ;
		RECT 18.710 25.360 18.890 25.695 ;
		LAYER VIA3 ;
		RECT 18.710 26.005 18.890 26.025 ;
		LAYER M2 ;
		RECT 18.710 39.280 18.890 39.615 ;
		LAYER M1 ;
		RECT 18.710 40.235 18.890 40.315 ;
		LAYER M2 ;
		RECT 18.710 40.255 18.890 40.295 ;
		LAYER M1 ;
		RECT 18.710 39.260 18.890 39.635 ;
		LAYER M3 ;
		RECT 18.710 39.925 18.890 39.945 ;
		LAYER M1 ;
		RECT 18.710 39.905 18.890 39.965 ;
		LAYER M3 ;
		RECT 18.710 40.255 18.890 40.295 ;
		LAYER M3 ;
		RECT 18.710 39.280 18.890 39.615 ;
		LAYER M3 ;
		RECT 18.710 40.935 18.890 41.290 ;
		LAYER VIA3 ;
		RECT 18.710 40.935 18.890 41.290 ;
		LAYER M1 ;
		RECT 18.710 38.265 18.890 38.325 ;
		LAYER M3 ;
		RECT 18.710 38.285 18.890 38.305 ;
		LAYER M2 ;
		RECT 18.710 38.285 18.890 38.305 ;
		LAYER VIA3 ;
		RECT 18.710 38.285 18.890 38.305 ;
		LAYER M2 ;
		RECT 18.710 40.605 18.890 40.625 ;
		LAYER M3 ;
		RECT 18.710 40.605 18.890 40.625 ;
		LAYER M1 ;
		RECT 18.710 40.585 18.890 40.645 ;
		LAYER M2 ;
		RECT 18.710 40.935 18.890 41.290 ;
		LAYER M2 ;
		RECT 18.710 38.615 18.890 38.970 ;
		LAYER M3 ;
		RECT 18.710 38.615 18.890 38.970 ;
		LAYER VIA3 ;
		RECT 18.710 38.615 18.890 38.970 ;
		LAYER M2 ;
		RECT 18.710 23.040 18.890 23.375 ;
		LAYER M1 ;
		RECT 18.710 23.020 18.890 23.395 ;
		LAYER M1 ;
		RECT 18.710 24.345 18.890 24.405 ;
		LAYER M1 ;
		RECT 18.710 23.665 18.890 23.725 ;
		LAYER VIA3 ;
		RECT 18.710 23.685 18.890 23.705 ;
		LAYER M3 ;
		RECT 18.710 24.365 18.890 24.385 ;
		LAYER M3 ;
		RECT 18.710 24.015 18.890 24.055 ;
		LAYER VIA3 ;
		RECT 18.710 24.015 18.890 24.055 ;
		LAYER M1 ;
		RECT 18.710 23.995 18.890 24.075 ;
		LAYER M2 ;
		RECT 18.710 24.365 18.890 24.385 ;
		LAYER VIA3 ;
		RECT 18.710 24.365 18.890 24.385 ;
		LAYER M3 ;
		RECT 18.710 12.415 18.890 12.455 ;
		LAYER M3 ;
		RECT 18.710 12.085 18.890 12.105 ;
		LAYER VIA3 ;
		RECT 18.710 12.085 18.890 12.105 ;
		LAYER M2 ;
		RECT 18.710 12.085 18.890 12.105 ;
		LAYER M3 ;
		RECT 18.710 7.445 18.890 7.465 ;
		LAYER VIA3 ;
		RECT 18.710 7.445 18.890 7.465 ;
		LAYER M3 ;
		RECT 18.710 6.135 18.890 6.490 ;
		LAYER M2 ;
		RECT 18.710 6.800 18.890 7.135 ;
		LAYER VIA3 ;
		RECT 18.710 6.135 18.890 6.490 ;
		LAYER M1 ;
		RECT 18.710 8.105 18.890 8.165 ;
		LAYER M2 ;
		RECT 18.710 5.805 18.890 5.825 ;
		LAYER M3 ;
		RECT 18.710 5.805 18.890 5.825 ;
		LAYER VIA3 ;
		RECT 18.710 5.805 18.890 5.825 ;
		LAYER M1 ;
		RECT 18.710 5.785 18.890 5.845 ;
		LAYER VIA3 ;
		RECT 18.710 12.415 18.890 12.455 ;
		LAYER M1 ;
		RECT 18.710 10.425 18.890 10.485 ;
		LAYER M1 ;
		RECT 18.710 10.755 18.890 11.150 ;
		LAYER M1 ;
		RECT 18.710 12.065 18.890 12.125 ;
		LAYER M3 ;
		RECT 18.710 11.440 18.890 11.775 ;
		LAYER M2 ;
		RECT 18.710 11.440 18.890 11.775 ;
		LAYER M1 ;
		RECT 18.710 11.420 18.890 11.795 ;
		LAYER VIA3 ;
		RECT 18.710 10.775 18.890 11.130 ;
		LAYER M3 ;
		RECT 18.710 31.655 18.890 32.010 ;
		LAYER M1 ;
		RECT 18.710 31.635 18.890 32.030 ;
		LAYER M3 ;
		RECT 18.710 33.295 18.890 33.335 ;
		LAYER M2 ;
		RECT 18.710 37.605 18.890 37.625 ;
		LAYER M2 ;
		RECT 18.710 24.015 18.890 24.055 ;
		LAYER M3 ;
		RECT 18.710 47.565 18.890 47.585 ;
		LAYER VIA3 ;
		RECT 18.710 47.215 18.890 47.255 ;
		LAYER M3 ;
		RECT 18.710 46.240 18.890 46.575 ;
		LAYER M2 ;
		RECT 18.710 47.565 18.890 47.585 ;
		LAYER VIA3 ;
		RECT 18.710 47.565 18.890 47.585 ;
		LAYER M3 ;
		RECT 18.710 23.685 18.890 23.705 ;
		LAYER M2 ;
		RECT 18.710 47.895 18.890 48.250 ;
		LAYER M3 ;
		RECT 18.710 47.895 18.890 48.250 ;
		LAYER M1 ;
		RECT 18.710 13.740 18.890 14.115 ;
		LAYER M1 ;
		RECT 18.710 14.385 18.890 14.445 ;
		LAYER M1 ;
		RECT 18.710 49.185 18.890 49.245 ;
		LAYER M1 ;
		RECT 18.710 49.515 18.890 49.595 ;
		LAYER M1 ;
		RECT 18.710 49.865 18.890 49.925 ;
		LAYER M1 ;
		RECT 18.710 50.195 18.890 50.590 ;
		LAYER M1 ;
		RECT 18.710 31.305 18.890 31.365 ;
		LAYER VIA3 ;
		RECT 18.710 44.565 18.890 44.585 ;
		LAYER M2 ;
		RECT 18.710 42.925 18.890 42.945 ;
		LAYER M2 ;
		RECT 18.710 44.565 18.890 44.585 ;
		LAYER M1 ;
		RECT 18.710 42.905 18.890 42.965 ;
		LAYER VIA3 ;
		RECT 18.710 43.255 18.890 43.610 ;
		LAYER M2 ;
		RECT 18.710 49.205 18.890 49.225 ;
		LAYER M3 ;
		RECT 18.710 49.205 18.890 49.225 ;
		LAYER VIA3 ;
		RECT 18.710 49.205 18.890 49.225 ;
		LAYER VIA3 ;
		RECT 18.710 47.895 18.890 48.250 ;
		LAYER M3 ;
		RECT 18.710 48.560 18.890 48.895 ;
		LAYER VIA3 ;
		RECT 18.710 48.560 18.890 48.895 ;
		LAYER M3 ;
		RECT 18.710 130.205 18.890 130.225 ;
		LAYER M2 ;
		RECT 18.710 121.920 18.890 122.255 ;
		LAYER M1 ;
		RECT 18.710 121.900 18.890 122.275 ;
		LAYER VIA3 ;
		RECT 18.710 113.615 18.890 113.655 ;
		LAYER M1 ;
		RECT 18.710 97.705 18.890 97.765 ;
		LAYER M2 ;
		RECT 18.710 97.375 18.890 97.415 ;
		LAYER M3 ;
		RECT 18.710 111.295 18.890 111.335 ;
		LAYER VIA3 ;
		RECT 18.710 111.295 18.890 111.335 ;
		LAYER M3 ;
		RECT 18.710 113.615 18.890 113.655 ;
		LAYER M1 ;
		RECT 18.710 96.380 18.890 96.755 ;
		LAYER M3 ;
		RECT 18.710 95.405 18.890 95.425 ;
		LAYER M3 ;
		RECT 18.710 129.855 18.890 129.895 ;
		LAYER VIA3 ;
		RECT 18.710 129.855 18.890 129.895 ;
		LAYER M2 ;
		RECT 18.710 129.855 18.890 129.895 ;
		LAYER VIA3 ;
		RECT 18.710 123.245 18.890 123.265 ;
		LAYER M4 ;
		RECT 5.490 111.655 18.505 113.295 ;
		LAYER M4 ;
		RECT 5.490 109.335 18.505 110.975 ;
		LAYER M4 ;
		RECT 5.490 107.015 18.505 108.655 ;
		LAYER M4 ;
		RECT 5.490 104.695 18.505 106.335 ;
		LAYER M4 ;
		RECT 0.000 100.155 18.505 101.595 ;
		LAYER M4 ;
		RECT 0.000 109.435 18.505 110.875 ;
		LAYER M4 ;
		RECT 0.000 111.755 18.505 113.195 ;
		LAYER M4 ;
		RECT 0.000 109.335 3.610 110.975 ;
		LAYER M4 ;
		RECT 0.000 111.655 3.610 113.295 ;
		LAYER M4 ;
		RECT 5.490 100.055 18.505 101.695 ;
		LAYER M4 ;
		RECT 5.490 102.375 18.505 104.015 ;
		LAYER M4 ;
		RECT 0.000 102.475 18.505 103.915 ;
		LAYER M4 ;
		RECT 0.000 107.115 18.505 108.555 ;
		LAYER M4 ;
		RECT 0.000 104.795 18.505 106.235 ;
		LAYER M4 ;
		RECT 5.490 52.215 18.505 53.855 ;
		LAYER M4 ;
		RECT 0.000 52.315 18.505 53.755 ;
		LAYER M4 ;
		RECT 0.000 54.635 18.505 56.075 ;
		LAYER M4 ;
		RECT 0.000 54.535 3.610 56.175 ;
		LAYER M4 ;
		RECT 0.000 49.895 3.610 51.535 ;
		LAYER M4 ;
		RECT 0.000 47.575 3.610 49.215 ;
		LAYER M4 ;
		RECT 0.000 52.215 3.610 53.855 ;
		LAYER M4 ;
		RECT 5.490 49.895 18.505 51.535 ;
		LAYER M4 ;
		RECT 0.000 49.995 18.505 51.435 ;
		LAYER M4 ;
		RECT 0.000 47.675 18.505 49.115 ;
		LAYER M4 ;
		RECT 5.490 47.575 18.505 49.215 ;
		LAYER M4 ;
		RECT 0.000 76.750 3.610 78.835 ;
		LAYER M4 ;
		RECT 0.000 74.595 3.610 76.330 ;
		LAYER M4 ;
		RECT 0.000 73.225 3.610 74.175 ;
		LAYER M4 ;
		RECT 0.000 64.135 3.610 65.405 ;
		LAYER M4 ;
		RECT 0.000 71.205 3.610 72.805 ;
		LAYER M4 ;
		RECT 0.000 68.250 3.610 70.785 ;
		LAYER M4 ;
		RECT 0.000 79.175 3.610 80.815 ;
		LAYER M4 ;
		RECT 0.000 90.775 3.610 92.415 ;
		LAYER M4 ;
		RECT 0.000 56.855 3.610 58.495 ;
		LAYER M4 ;
		RECT 5.490 97.735 18.505 99.375 ;
		LAYER M4 ;
		RECT 0.000 97.835 18.505 99.275 ;
		LAYER M4 ;
		RECT 5.490 79.175 18.505 80.815 ;
		LAYER M4 ;
		RECT 0.000 76.850 18.505 78.785 ;
		LAYER M4 ;
		RECT 5.490 95.415 18.505 97.055 ;
		LAYER M4 ;
		RECT 0.000 97.735 3.610 99.375 ;
		LAYER M4 ;
		RECT 0.000 95.415 3.610 97.055 ;
		LAYER M4 ;
		RECT 0.000 74.695 18.505 76.230 ;
		LAYER M4 ;
		RECT 5.490 83.815 18.505 85.455 ;
		LAYER M4 ;
		RECT 0.000 83.915 18.505 85.355 ;
		LAYER M4 ;
		RECT 0.000 81.595 18.505 83.035 ;
		LAYER M4 ;
		RECT 5.490 81.495 18.505 83.135 ;
		LAYER M4 ;
		RECT 0.000 83.815 3.610 85.455 ;
		LAYER M4 ;
		RECT 0.000 81.495 3.610 83.135 ;
		LAYER M4 ;
		RECT 0.000 86.135 3.610 87.775 ;
		LAYER M4 ;
		RECT 5.490 86.135 18.505 87.775 ;
		LAYER M4 ;
		RECT 0.000 88.555 18.505 89.995 ;
		LAYER M4 ;
		RECT 5.490 88.455 18.505 90.095 ;
		LAYER M4 ;
		RECT 0.000 88.455 3.610 90.095 ;
		LAYER M4 ;
		RECT 0.000 86.235 18.505 87.675 ;
		LAYER M4 ;
		RECT 5.490 90.775 18.505 92.415 ;
		LAYER M4 ;
		RECT 0.000 90.875 18.505 92.315 ;
		LAYER M4 ;
		RECT 0.000 79.275 18.505 80.715 ;
		LAYER M4 ;
		RECT 0.000 93.095 3.610 94.735 ;
		LAYER M4 ;
		RECT 5.490 93.095 18.505 94.735 ;
		LAYER M4 ;
		RECT 0.000 93.195 18.505 94.635 ;
		LAYER M4 ;
		RECT 0.000 95.515 18.505 96.955 ;
		LAYER M4 ;
		RECT 5.490 76.750 16.685 78.160 ;
		LAYER M4 ;
		RECT 5.490 64.135 18.555 65.405 ;
		LAYER M4 ;
		RECT 5.490 62.555 18.555 63.715 ;
		LAYER M4 ;
		RECT 5.490 74.595 18.555 76.330 ;
		LAYER M4 ;
		RECT 5.490 73.225 18.555 74.175 ;
		LAYER M4 ;
		RECT 5.490 71.205 18.555 72.805 ;
		LAYER M4 ;
		RECT 5.490 68.250 18.555 70.785 ;
		LAYER M4 ;
		RECT 5.490 65.825 18.555 67.830 ;
		LAYER M4 ;
		RECT 16.685 76.750 18.555 77.930 ;
		LAYER M4 ;
		RECT 16.685 61.670 18.555 62.135 ;
		LAYER M4 ;
		RECT 0.000 73.325 18.505 74.075 ;
		LAYER M4 ;
		RECT 0.000 68.350 18.505 70.685 ;
		LAYER M4 ;
		RECT 0.000 71.305 18.505 72.705 ;
		LAYER M4 ;
		RECT 0.000 62.555 3.610 63.715 ;
		LAYER M4 ;
		RECT 5.490 61.520 16.685 62.135 ;
		LAYER M4 ;
		RECT 0.000 58.885 18.505 62.035 ;
		LAYER M4 ;
		RECT 5.490 56.855 18.505 58.495 ;
		LAYER M4 ;
		RECT 0.000 61.670 3.610 62.135 ;
		LAYER M4 ;
		RECT 0.000 65.825 3.610 67.830 ;
		LAYER M4 ;
		RECT 0.000 65.925 18.555 67.730 ;
		LAYER M4 ;
		RECT 0.000 64.235 18.555 65.305 ;
		LAYER M4 ;
		RECT 0.000 62.655 18.555 63.615 ;
		LAYER M3 ;
		RECT 18.710 35.285 18.890 35.305 ;
		LAYER M2 ;
		RECT 18.710 35.285 18.890 35.305 ;
		LAYER M2 ;
		RECT 18.710 34.640 18.890 34.975 ;
		LAYER M3 ;
		RECT 18.710 34.640 18.890 34.975 ;
		LAYER M1 ;
		RECT 18.710 37.585 18.890 37.645 ;
		LAYER M4 ;
		RECT 5.490 35.975 18.505 37.615 ;
		LAYER M4 ;
		RECT 0.000 36.075 18.505 37.515 ;
		LAYER M4 ;
		RECT 0.000 38.395 18.505 39.835 ;
		LAYER M4 ;
		RECT 0.000 35.975 3.610 37.615 ;
		LAYER M4 ;
		RECT 0.000 38.295 3.610 39.935 ;
		LAYER M4 ;
		RECT 5.490 45.255 18.505 46.895 ;
		LAYER M4 ;
		RECT 0.000 45.355 18.505 46.795 ;
		LAYER M4 ;
		RECT 0.000 43.035 18.505 44.475 ;
		LAYER M4 ;
		RECT 5.490 42.935 18.505 44.575 ;
		LAYER M4 ;
		RECT 0.000 42.935 3.610 44.575 ;
		LAYER M4 ;
		RECT 5.490 33.655 18.505 35.295 ;
		LAYER M4 ;
		RECT 0.000 33.755 18.505 35.195 ;
		LAYER M4 ;
		RECT 0.000 33.655 3.610 35.295 ;
		LAYER M4 ;
		RECT 5.490 31.335 18.505 32.975 ;
		LAYER M4 ;
		RECT 0.000 31.335 3.610 32.975 ;
		LAYER M4 ;
		RECT 0.000 31.435 18.505 32.875 ;
		LAYER M4 ;
		RECT 0.000 29.015 3.610 30.655 ;
		LAYER M4 ;
		RECT 5.490 29.015 18.505 30.655 ;
		LAYER M4 ;
		RECT 5.490 26.695 18.505 28.335 ;
		LAYER M4 ;
		RECT 0.000 26.795 18.505 28.235 ;
		LAYER M4 ;
		RECT 0.000 26.695 3.610 28.335 ;
		LAYER M4 ;
		RECT 0.000 29.115 18.505 30.555 ;
		LAYER M4 ;
		RECT 0.000 45.255 3.610 46.895 ;
		LAYER M4 ;
		RECT 0.000 40.615 3.610 42.255 ;
		LAYER M4 ;
		RECT 0.000 40.715 18.505 42.155 ;
		LAYER M4 ;
		RECT 5.490 40.615 18.505 42.255 ;
		LAYER M4 ;
		RECT 0.000 127.895 3.610 129.535 ;
		LAYER M4 ;
		RECT 0.000 100.055 3.610 101.695 ;
		LAYER M4 ;
		RECT 0.000 102.375 3.610 104.015 ;
		LAYER M4 ;
		RECT 0.000 104.695 3.610 106.335 ;
		LAYER M4 ;
		RECT 0.000 123.255 3.610 124.895 ;
		LAYER M4 ;
		RECT 0.000 120.935 3.610 122.575 ;
		LAYER M4 ;
		RECT 0.000 113.975 3.610 115.615 ;
		LAYER M4 ;
		RECT 0.000 107.015 3.610 108.655 ;
		LAYER M4 ;
		RECT 5.490 113.975 18.505 115.615 ;
		LAYER M4 ;
		RECT 5.490 116.295 18.505 117.935 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 18.710 137.670 ;
		LAYER M4 ;
		RECT 0.000 0.000 18.505 0.785 ;
		LAYER M4 ;
		RECT 5.490 24.375 18.505 26.015 ;
		LAYER M4 ;
		RECT 5.490 1.175 18.505 2.815 ;
		LAYER M4 ;
		RECT 5.490 3.495 18.505 5.135 ;
		LAYER M4 ;
		RECT 0.000 1.175 3.610 2.815 ;
		LAYER M4 ;
		RECT 0.000 1.275 18.505 2.715 ;
		LAYER M4 ;
		RECT 5.490 15.095 18.505 16.735 ;
		LAYER M4 ;
		RECT 5.490 12.775 18.505 14.415 ;
		LAYER M4 ;
		RECT 5.490 10.455 18.505 12.095 ;
		LAYER M4 ;
		RECT 5.490 8.135 18.505 9.775 ;
		LAYER M4 ;
		RECT 5.490 19.735 18.505 21.375 ;
		LAYER M4 ;
		RECT 5.490 17.415 18.505 19.055 ;
		LAYER M4 ;
		RECT 0.000 17.515 18.505 18.955 ;
		LAYER M4 ;
		RECT 0.000 15.195 18.505 16.635 ;
		LAYER M4 ;
		RECT 0.000 22.055 3.610 23.695 ;
		LAYER M4 ;
		RECT 0.000 22.155 18.505 23.595 ;
		LAYER M4 ;
		RECT 0.000 24.475 18.505 25.915 ;
		LAYER M4 ;
		RECT 5.490 22.055 18.505 23.695 ;
		LAYER M4 ;
		RECT 0.000 24.375 3.610 26.015 ;
		LAYER M4 ;
		RECT 18.555 0.000 18.890 137.670 ;
		LAYER M4 ;
		RECT 18.505 0.000 18.555 62.035 ;
		LAYER M3 ;
		RECT 0.000 0.000 18.710 137.670 ;
		LAYER M1 ;
		RECT 0.000 0.000 18.710 137.670 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 18.890 137.670 ;
		LAYER M4 ;
		RECT 5.490 123.255 18.505 124.895 ;
		LAYER M4 ;
		RECT 0.000 123.355 18.505 124.795 ;
		LAYER M4 ;
		RECT 5.490 125.575 18.505 127.215 ;
		LAYER M4 ;
		RECT 0.000 127.995 18.505 129.435 ;
		LAYER M4 ;
		RECT 5.490 132.535 18.505 134.175 ;
		LAYER M4 ;
		RECT 0.000 132.635 18.505 134.075 ;
		LAYER M4 ;
		RECT 0.000 134.955 18.505 136.395 ;
		LAYER M4 ;
		RECT 5.490 134.855 18.505 136.495 ;
		LAYER M4 ;
		RECT 0.000 130.215 3.610 131.855 ;
		LAYER M4 ;
		RECT 5.490 130.215 18.505 131.855 ;
		LAYER M4 ;
		RECT 0.000 130.315 18.505 131.755 ;
		LAYER M4 ;
		RECT 5.490 120.935 18.505 122.575 ;
		LAYER M2 ;
		RECT 0.000 0.000 18.710 137.670 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 18.890 137.670 ;
		LAYER M4 ;
		RECT 5.490 54.535 18.505 56.175 ;
		LAYER M4 ;
		RECT 0.000 56.955 18.505 58.395 ;
		LAYER M4 ;
		RECT 5.490 38.295 18.505 39.935 ;
		LAYER M4 ;
		RECT 5.490 127.895 18.505 129.535 ;
		LAYER M4 ;
		RECT 0.000 116.395 18.505 117.835 ;
		LAYER M4 ;
		RECT 0.000 114.075 18.505 115.515 ;
		LAYER M4 ;
		RECT 0.000 134.855 3.610 136.495 ;
		LAYER M4 ;
		RECT 0.000 132.535 3.610 134.175 ;
		LAYER M4 ;
		RECT 0.000 136.885 18.505 137.670 ;
		LAYER M4 ;
		RECT 0.000 118.615 3.610 120.255 ;
		LAYER M4 ;
		RECT 0.000 116.295 3.610 117.935 ;
		LAYER M4 ;
		RECT 0.000 125.575 3.610 127.215 ;
		LAYER M4 ;
		RECT 0.000 125.675 18.505 127.115 ;
		LAYER M4 ;
		RECT 0.000 121.035 18.505 122.475 ;
		LAYER M4 ;
		RECT 0.000 118.715 18.505 120.155 ;
		LAYER M4 ;
		RECT 5.490 118.615 18.505 120.255 ;
		LAYER M4 ;
		RECT 0.000 19.735 3.610 21.375 ;
		LAYER M4 ;
		RECT 0.000 15.095 3.610 16.735 ;
		LAYER M4 ;
		RECT 0.000 17.415 3.610 19.055 ;
		LAYER M4 ;
		RECT 0.000 19.835 18.505 21.275 ;
		LAYER M4 ;
		RECT 0.000 10.455 3.610 12.095 ;
		LAYER M4 ;
		RECT 0.000 8.135 3.610 9.775 ;
		LAYER M4 ;
		RECT 0.000 5.815 3.610 7.455 ;
		LAYER M4 ;
		RECT 0.000 12.775 3.610 14.415 ;
		LAYER M4 ;
		RECT 5.490 5.815 18.505 7.455 ;
		LAYER M4 ;
		RECT 0.000 5.915 18.505 7.355 ;
		LAYER M4 ;
		RECT 0.000 8.235 18.505 9.675 ;
		LAYER M4 ;
		RECT 0.000 10.555 18.505 11.995 ;
		LAYER M4 ;
		RECT 0.000 3.495 3.610 5.135 ;
		LAYER M4 ;
		RECT 0.000 3.595 18.505 5.035 ;
		LAYER M4 ;
		RECT 0.000 12.875 18.505 14.315 ;
	END
	# End of OBS

END TS1N28HPCPUHDHVTB32X50M4SWBSO

END LIBRARY
